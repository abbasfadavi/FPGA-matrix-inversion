LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY SinglePortRAM_generic IS
  GENERIC( AddrWidth                      : integer := 1;
           DataWidth                      : integer := 1
           );
  PORT( clk                               :   IN    std_logic;
        din_re                            :   IN    std_logic_vector(DataWidth - 1 DOWNTO 0);
        din_im                            :   IN    std_logic_vector(DataWidth - 1 DOWNTO 0);
        addr                              :   IN    std_logic_vector(AddrWidth - 1 DOWNTO 0);
        we                                :   IN    std_logic;
        dout_re                           :   OUT   std_logic_vector(DataWidth - 1 DOWNTO 0);
        dout_im                           :   OUT   std_logic_vector(DataWidth - 1 DOWNTO 0)
        );
END SinglePortRAM_generic;


ARCHITECTURE rtl OF SinglePortRAM_generic IS

  -- Local Type Definitions
  TYPE ram_type IS ARRAY (2**AddrWidth - 1 DOWNTO 0) of std_logic_vector(DataWidth*2 - 1 DOWNTO 0);

  -- Signals
  SIGNAL ram                              : ram_type;
  SIGNAL data_int                         : std_logic_vector(DataWidth*2 - 1 DOWNTO 0);
  SIGNAL addr_unsigned                    : unsigned(AddrWidth - 1 DOWNTO 0);

BEGIN
  addr_unsigned <= unsigned(addr);

  SinglePortRAM_generic_process: PROCESS (clk)
  BEGIN
    IF clk'event AND clk = '1' THEN
      IF we = '1' THEN
        ram(to_integer(addr_unsigned)) <= din_re & din_im;
        data_int <= din_re & din_im;
      ELSE
        data_int <= ram(to_integer(addr_unsigned));
      END IF;
    END IF;
  END PROCESS SinglePortRAM_generic_process;

  dout_re <= data_int(DataWidth*2-1 DOWNTO DataWidth);
  dout_im <= data_int(DataWidth-1 DOWNTO 0);

END rtl;

