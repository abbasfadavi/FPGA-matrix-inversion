LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.my_inverse_pac.ALL;

ENTITY nfp_sub_single IS
  PORT( clk                               :   IN    std_logic;
        reset_x                           :   IN    std_logic;
        enb                               :   IN    std_logic;
        nfp_in1                           :   IN    std_logic_vector(31 DOWNTO 0);
        nfp_in2                           :   IN    std_logic_vector(31 DOWNTO 0);
        nfp_out                           :   OUT   std_logic_vector(31 DOWNTO 0)
        );
END nfp_sub_single;


ARCHITECTURE rtl OF nfp_sub_single IS

  -- Signals
  SIGNAL nfp_in1_unsigned                 : unsigned(31 DOWNTO 0);
  SIGNAL AS                               : std_logic;
  SIGNAL AE                               : unsigned(7 DOWNTO 0);
  SIGNAL AM                               : unsigned(22 DOWNTO 0);
  SIGNAL Delay1_out1                      : unsigned(7 DOWNTO 0);
  SIGNAL nfp_in2_unsigned                 : unsigned(31 DOWNTO 0);
  SIGNAL BS                               : std_logic;
  SIGNAL BE                               : unsigned(7 DOWNTO 0);
  SIGNAL BM                               : unsigned(22 DOWNTO 0);
  SIGNAL Delay4_out1                      : unsigned(7 DOWNTO 0);
  SIGNAL Relational_Operator1_relop1      : std_logic;
  SIGNAL Delay2_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL Delay5_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL Relational_Operator_relop1       : std_logic;
  SIGNAL bitconcat_aExponent_aMantissa_relop1 : std_logic;
  SIGNAL Logical_Operator_out1            : std_logic;
  SIGNAL Logical_Operator1_out1           : std_logic;
  SIGNAL if_bitconcat_aExponent_aMantiss_out1 : unsigned(7 DOWNTO 0);
  SIGNAL aExponent_cfType_Exponent_I_out1 : std_logic;
  SIGNAL Delay11_out1                     : std_logic;
  SIGNAL Delay42_out1                     : std_logic;
  SIGNAL Delay18_reg_rsvd                 : std_logic_vector(0 TO 1);
  SIGNAL Delay18_reg_next                 : std_logic_vector(0 TO 1);
  SIGNAL Delay18_out1                     : std_logic;
  SIGNAL Exponent_0_out1                  : std_logic;
  SIGNAL C_out1                           : unsigned(7 DOWNTO 0);
  SIGNAL if_Exponent_0_out1               : unsigned(7 DOWNTO 0);
  SIGNAL Delay_out1                       : unsigned(7 DOWNTO 0);
  SIGNAL Delay4_out1_1                    : unsigned(7 DOWNTO 0);
  SIGNAL Delay2_out1_1                    : unsigned(7 DOWNTO 0);
  SIGNAL exp_norm_cfType_Exponent_In_out1 : std_logic;
  SIGNAL alphaExponent_0_cfType_Exp_out1  : std_logic;
  SIGNAL alpha1_out1                      : unsigned(2 DOWNTO 0);
  SIGNAL alpha0_out1                      : unsigned(2 DOWNTO 0);
  SIGNAL if_Exponent_0_cfType_Exp_out1    : unsigned(2 DOWNTO 0);
  SIGNAL if_bitconcat_aExponent_aMantiss_1_ou_1 : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Concat_out1                  : unsigned(25 DOWNTO 0);
  SIGNAL alpha0_1_out1                    : unsigned(1 DOWNTO 0);
  SIGNAL Bit_Concat1_out1                 : unsigned(27 DOWNTO 0);
  SIGNAL Data_Type_Conversion_out1        : signed(27 DOWNTO 0);
  SIGNAL Delay2_out1_2                    : signed(27 DOWNTO 0);
  SIGNAL Delay5_out1_1                    : signed(27 DOWNTO 0);
  SIGNAL Delay3_out1                      : std_logic;
  SIGNAL Logical_Operator_out1_1          : std_logic;
  SIGNAL Delay_out1_1                     : std_logic;
  SIGNAL if_bitconcat_aExponent_aMantiss_2_ou_1 : std_logic;
  SIGNAL if_bitconcat_aExponent_aMantiss_5_ou_1 : std_logic;
  SIGNAL bitxor_out1                      : std_logic;
  SIGNAL Delay10_out1                     : std_logic;
  SIGNAL if_bitconcat_aExponent_aMantiss_3_ou_1 : unsigned(7 DOWNTO 0);
  SIGNAL exp_b_cfType_Exponent_Inf_o_out1 : std_logic;
  SIGNAL Exponent_0_out1_1                : std_logic;
  SIGNAL alphaExponent_0_cfType_Exp_out1_1 : std_logic;
  SIGNAL alpha1_out1_1                    : unsigned(2 DOWNTO 0);
  SIGNAL alpha0_out1_1                    : unsigned(2 DOWNTO 0);
  SIGNAL if_Exponent_0_cfType_Exp_out1_1  : unsigned(2 DOWNTO 0);
  SIGNAL if_bitconcat_aExponent_aMantiss_4_ou_1 : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Concat_out1_1                : unsigned(25 DOWNTO 0);
  SIGNAL alpha0_1_out1_1                  : unsigned(1 DOWNTO 0);
  SIGNAL Bit_Concat1_out1_1               : unsigned(27 DOWNTO 0);
  SIGNAL Data_Type_Conversion_out1_1      : signed(27 DOWNTO 0);
  SIGNAL Delay1_out1_1                    : signed(27 DOWNTO 0);
  SIGNAL alphamant_b_ext_in0              : signed(28 DOWNTO 0);
  SIGNAL alphamant_b_ext_out1             : signed(27 DOWNTO 0);
  SIGNAL if_opp_Sign_out1                 : signed(27 DOWNTO 0);
  SIGNAL C_out1_1                         : unsigned(7 DOWNTO 0);
  SIGNAL if_Exponent_0_out1_1             : unsigned(7 DOWNTO 0);
  SIGNAL Delay_out1_2                     : unsigned(7 DOWNTO 0);
  SIGNAL storedInteger_exp_a_cor_sto_sub_cast : signed(31 DOWNTO 0);
  SIGNAL storedInteger_exp_a_cor_sto_sub_cast_1 : signed(31 DOWNTO 0);
  SIGNAL storedInteger_exp_a_cor_sto_out1 : signed(31 DOWNTO 0);
  SIGNAL Bit_Slice2_out1                  : unsigned(2 DOWNTO 0);
  SIGNAL Compare_To_Zero_out1             : std_logic;
  SIGNAL Constant_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Bit_Slice_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL if_opp_Sign_1_out1               : unsigned(4 DOWNTO 0);
  SIGNAL bitsra_mant_b_ext_shift_lengt_out1 : signed(27 DOWNTO 0);
  SIGNAL Delay1_out1_2                    : signed(27 DOWNTO 0);
  SIGNAL mant_a_ext_mant_b_shifted_add_temp : signed(31 DOWNTO 0);
  SIGNAL mant_a_ext_mant_b_shifted_out1   : unsigned(26 DOWNTO 0);
  SIGNAL BitSlice_out1                    : std_logic;
  SIGNAL Delay3_out1_1                    : std_logic;
  SIGNAL Logical_Operator_out1_2          : std_logic;
  SIGNAL Delay13_out1                     : std_logic;
  SIGNAL Delay1_out1_3                    : unsigned(26 DOWNTO 0);
  SIGNAL BitSlice3_out1                   : unsigned(25 DOWNTO 0);
  SIGNAL Bit_Slice5_out1                  : std_logic;
  SIGNAL Bit_Slice3_out1                  : std_logic;
  SIGNAL Logical_Operator1_out1_1         : std_logic;
  SIGNAL Bit_Slice2_out1_1                : unsigned(7 DOWNTO 0);
  SIGNAL Bit_Slice16_out1                 : std_logic;
  SIGNAL Bit_Slice15_out1                 : std_logic;
  SIGNAL Logical_Operator5_out1           : std_logic;
  SIGNAL Bit_Slice14_out1                 : std_logic;
  SIGNAL Bit_Slice13_out1                 : std_logic;
  SIGNAL Logical_Operator7_out1           : std_logic;
  SIGNAL Logical_Operator6_out1           : std_logic;
  SIGNAL Bit_Slice12_out1                 : std_logic;
  SIGNAL Bit_Slice11_out1                 : std_logic;
  SIGNAL Logical_Operator4_out1           : std_logic;
  SIGNAL Bit_Slice10_out1                 : std_logic;
  SIGNAL Bit_Slice9_out1                  : std_logic;
  SIGNAL Logical_Operator14_out1          : std_logic;
  SIGNAL Logical_Operator13_out1          : std_logic;
  SIGNAL Logical_Operator12_out1          : std_logic;
  SIGNAL Bit_Slice1_out1                  : unsigned(7 DOWNTO 0);
  SIGNAL Bit_Slice16_out1_1               : std_logic;
  SIGNAL Bit_Slice15_out1_1               : std_logic;
  SIGNAL Logical_Operator5_out1_1         : std_logic;
  SIGNAL Bit_Slice14_out1_1               : std_logic;
  SIGNAL Bit_Slice13_out1_1               : std_logic;
  SIGNAL Logical_Operator7_out1_1         : std_logic;
  SIGNAL Logical_Operator6_out1_1         : std_logic;
  SIGNAL Bit_Slice12_out1_1               : std_logic;
  SIGNAL Bit_Slice11_out1_1               : std_logic;
  SIGNAL Logical_Operator4_out1_1         : std_logic;
  SIGNAL Bit_Slice10_out1_1               : std_logic;
  SIGNAL Bit_Slice9_out1_1                : std_logic;
  SIGNAL Logical_Operator14_out1_1        : std_logic;
  SIGNAL Logical_Operator13_out1_1        : std_logic;
  SIGNAL Bit_Slice4_out1                  : unsigned(7 DOWNTO 0);
  SIGNAL Bit_Slice8_out1                  : std_logic;
  SIGNAL Bit_Slice7_out1                  : std_logic;
  SIGNAL Logical_Operator1_out1_2         : std_logic;
  SIGNAL Bit_Slice6_out1                  : std_logic;
  SIGNAL Bit_Slice5_out1_1                : std_logic;
  SIGNAL Logical_Operator3_out1           : std_logic;
  SIGNAL Bit_Slice3_out1_1                : std_logic;
  SIGNAL Bit_Slice2_out1_2                : std_logic;
  SIGNAL Bit_Slice1_out1_1                : std_logic;
  SIGNAL Bit_Slice_out1_1                 : std_logic;
  SIGNAL Constant_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant1_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch_out1                      : unsigned(4 DOWNTO 0);
  SIGNAL Logical_Operator_out1_3          : std_logic;
  SIGNAL Constant2_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch1_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant3_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch2_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant4_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Logical_Operator2_out1           : std_logic;
  SIGNAL Switch3_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Switch4_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant5_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch5_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant6_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch6_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant7_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch7_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Constant8_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch8_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Logical_Operator12_out1_1        : std_logic;
  SIGNAL Switch9_out1                     : unsigned(4 DOWNTO 0);
  SIGNAL Switch10_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant9_out1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch11_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant10_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch12_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant11_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch14_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant12_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch15_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Switch16_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant13_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch17_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant14_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch18_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant15_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch19_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant16_out1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch20_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Switch21_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Logical_Operator_out1_4          : std_logic;
  SIGNAL Switch13_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Switch33_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Constant9_out1_1                 : unsigned(4 DOWNTO 0);
  SIGNAL Switch11_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant10_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch12_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant11_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch14_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant12_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch15_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch16_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant13_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch17_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant14_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch18_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant15_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch19_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant16_out1_1                : unsigned(4 DOWNTO 0);
  SIGNAL Switch20_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch21_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Switch13_out1_1                  : unsigned(4 DOWNTO 0);
  SIGNAL Constant1_out1_1                 : unsigned(4 DOWNTO 0);
  SIGNAL Switch3_out1_1                   : unsigned(4 DOWNTO 0);
  SIGNAL Constant2_out1_1                 : unsigned(4 DOWNTO 0);
  SIGNAL Switch2_out1_1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch1_out1_1                   : unsigned(4 DOWNTO 0);
  SIGNAL Switch34_out1                    : unsigned(4 DOWNTO 0);
  SIGNAL Delay_out1_3                     : unsigned(4 DOWNTO 0);
  SIGNAL Bit_Slice_out1_2                 : unsigned(4 DOWNTO 0);
  SIGNAL shift_length_exp_a_cor_relop1    : std_logic;
  SIGNAL Bit_Slice1_out1_2                : unsigned(2 DOWNTO 0);
  SIGNAL Compare_To_Zero_out1_1           : std_logic;
  SIGNAL Logical_Operator1_out1_3         : std_logic;
  SIGNAL C1_out1                          : unsigned(7 DOWNTO 0);
  SIGNAL exp_a_cor_1_out1                 : unsigned(4 DOWNTO 0);
  SIGNAL if_shift_length_exp_a_cor_1_out1 : unsigned(4 DOWNTO 0);
  SIGNAL bitsll_Sum_shift_length_out1     : unsigned(26 DOWNTO 0);
  SIGNAL bitsrl_Sum_1_out1                : unsigned(26 DOWNTO 0);
  SIGNAL if_bitget_Sum_Sum_WordLength_out1 : unsigned(26 DOWNTO 0);
  SIGNAL Delay15_out1                     : unsigned(26 DOWNTO 0);
  SIGNAL C5_out1                          : unsigned(26 DOWNTO 0);
  SIGNAL if_exp_norm_cfType_Exponent_I_out1 : unsigned(26 DOWNTO 0);
  SIGNAL BitSlice6_out1                   : unsigned(23 DOWNTO 0);
  SIGNAL BitSlice5_out1                   : std_logic;
  SIGNAL Bit_Slice13_out1_2               : std_logic;
  SIGNAL Bit_Slice12_out1_2               : std_logic;
  SIGNAL Bit_Slice10_out1_2               : std_logic;
  SIGNAL Bit_Slice11_out1_2               : std_logic;
  SIGNAL Bit_Slice14_out1_2               : std_logic;
  SIGNAL Bit_Slice7_out1_1                : unsigned(2 DOWNTO 0);
  SIGNAL Constant1_out1_2                 : std_logic;
  SIGNAL Bit_Concat_out1_2                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_3                 : std_logic;
  SIGNAL Data_Type_Conversion_out1_2      : std_logic;
  SIGNAL Bit_Slice1_out1_3                : std_logic;
  SIGNAL Logical_Operator_out1_5          : std_logic;
  SIGNAL Switch6_out1_1                   : std_logic;
  SIGNAL Bit_Slice2_out1_3                : std_logic;
  SIGNAL Logical_Operator1_out1_4         : std_logic;
  SIGNAL Bit_Slice3_out1_2                : std_logic;
  SIGNAL Logical_Operator2_out1_1         : std_logic;
  SIGNAL Switch7_out1_1                   : std_logic;
  SIGNAL Switch3_out1_2                   : std_logic;
  SIGNAL Bit_Slice8_out1_1                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_4                 : std_logic;
  SIGNAL Logical_Operator3_out1_1         : std_logic;
  SIGNAL Bit_Slice1_out1_4                : std_logic;
  SIGNAL Logical_Operator_out1_6          : std_logic;
  SIGNAL Switch6_out1_2                   : std_logic;
  SIGNAL Bit_Slice2_out1_4                : std_logic;
  SIGNAL Logical_Operator1_out1_5         : std_logic;
  SIGNAL Bit_Slice3_out1_3                : std_logic;
  SIGNAL Logical_Operator2_out1_2         : std_logic;
  SIGNAL Switch7_out1_2                   : std_logic;
  SIGNAL Switch3_out1_3                   : std_logic;
  SIGNAL Switch6_out1_3                   : std_logic;
  SIGNAL Bit_Slice9_out1_2                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_5                 : std_logic;
  SIGNAL Logical_Operator3_out1_2         : std_logic;
  SIGNAL Bit_Slice1_out1_5                : std_logic;
  SIGNAL Logical_Operator_out1_7          : std_logic;
  SIGNAL Switch6_out1_4                   : std_logic;
  SIGNAL Bit_Slice2_out1_5                : std_logic;
  SIGNAL Logical_Operator1_out1_6         : std_logic;
  SIGNAL Bit_Slice3_out1_4                : std_logic;
  SIGNAL Logical_Operator2_out1_3         : std_logic;
  SIGNAL Switch7_out1_3                   : std_logic;
  SIGNAL Switch3_out1_4                   : std_logic;
  SIGNAL Bit_Slice3_out1_5                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_6                 : std_logic;
  SIGNAL Logical_Operator3_out1_3         : std_logic;
  SIGNAL Bit_Slice1_out1_6                : std_logic;
  SIGNAL Logical_Operator_out1_8          : std_logic;
  SIGNAL Switch6_out1_5                   : std_logic;
  SIGNAL Bit_Slice2_out1_6                : std_logic;
  SIGNAL Logical_Operator1_out1_7         : std_logic;
  SIGNAL Bit_Slice3_out1_6                : std_logic;
  SIGNAL Logical_Operator2_out1_4         : std_logic;
  SIGNAL Switch7_out1_4                   : std_logic;
  SIGNAL Switch3_out1_5                   : std_logic;
  SIGNAL Switch7_out1_5                   : std_logic;
  SIGNAL Switch3_out1_6                   : std_logic;
  SIGNAL Bit_Slice4_out1_1                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_7                 : std_logic;
  SIGNAL Logical_Operator3_out1_4         : std_logic;
  SIGNAL Bit_Slice1_out1_7                : std_logic;
  SIGNAL Logical_Operator_out1_9          : std_logic;
  SIGNAL Switch6_out1_6                   : std_logic;
  SIGNAL Bit_Slice2_out1_7                : std_logic;
  SIGNAL Logical_Operator1_out1_8         : std_logic;
  SIGNAL Bit_Slice3_out1_7                : std_logic;
  SIGNAL Logical_Operator2_out1_5         : std_logic;
  SIGNAL Switch7_out1_6                   : std_logic;
  SIGNAL Switch3_out1_7                   : std_logic;
  SIGNAL Bit_Slice5_out1_2                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_8                 : std_logic;
  SIGNAL Logical_Operator3_out1_5         : std_logic;
  SIGNAL Bit_Slice1_out1_8                : std_logic;
  SIGNAL Logical_Operator_out1_10         : std_logic;
  SIGNAL Switch6_out1_7                   : std_logic;
  SIGNAL Bit_Slice2_out1_8                : std_logic;
  SIGNAL Logical_Operator1_out1_9         : std_logic;
  SIGNAL Bit_Slice3_out1_8                : std_logic;
  SIGNAL Logical_Operator2_out1_6         : std_logic;
  SIGNAL Switch7_out1_7                   : std_logic;
  SIGNAL Switch3_out1_8                   : std_logic;
  SIGNAL Switch6_out1_8                   : std_logic;
  SIGNAL Bit_Slice6_out1_1                : unsigned(3 DOWNTO 0);
  SIGNAL Bit_Slice_out1_9                 : std_logic;
  SIGNAL Logical_Operator3_out1_6         : std_logic;
  SIGNAL Bit_Slice1_out1_9                : std_logic;
  SIGNAL Logical_Operator_out1_11         : std_logic;
  SIGNAL Switch6_out1_9                   : std_logic;
  SIGNAL Bit_Slice2_out1_9                : std_logic;
  SIGNAL Logical_Operator1_out1_10        : std_logic;
  SIGNAL Bit_Slice3_out1_9                : std_logic;
  SIGNAL Logical_Operator2_out1_7         : std_logic;
  SIGNAL Switch7_out1_8                   : std_logic;
  SIGNAL Switch3_out1_9                   : std_logic;
  SIGNAL Bit_Slice1_out1_10               : std_logic;
  SIGNAL Logical_Operator_out1_12         : std_logic;
  SIGNAL Logical_Operator1_out1_11        : std_logic;
  SIGNAL Switch7_out1_9                   : std_logic;
  SIGNAL Switch3_out1_10                  : std_logic;
  SIGNAL Switch2_out1_2                   : std_logic;
  SIGNAL Delay_out1_4                     : std_logic;
  SIGNAL Delay12_out1                     : std_logic;
  SIGNAL BitSlice1_out1                   : std_logic;
  SIGNAL sticky_bitget_Sum_1_out1         : std_logic;
  SIGNAL Delay4_out1_2                    : std_logic;
  SIGNAL if_bitget_Sum_Sum_WordLength_2_out1 : std_logic;
  SIGNAL BitSlice_out1_1                  : std_logic;
  SIGNAL BitSlice1_out1_1                 : std_logic;
  SIGNAL Delay19_out1                     : std_logic;
  SIGNAL sticky_bitget_Sum_1_out1_1       : std_logic;
  SIGNAL alphabitget_Mant_tmp_2_0_out1    : std_logic;
  SIGNAL alphabitget_Mant_tmp_1_0_out1    : std_logic;
  SIGNAL alpha0_out1_2                    : std_logic;
  SIGNAL BitSlice4_out1                   : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Concat_out1_3                : unsigned(23 DOWNTO 0);
  SIGNAL cast_2_like_Mant_tmp_out1        : unsigned(23 DOWNTO 0);
  SIGNAL Mant_tmp_cast_2_like_Man_out1    : unsigned(23 DOWNTO 0);
  SIGNAL if_bitget_Mant_tmp_1_0_out1      : unsigned(23 DOWNTO 0);
  SIGNAL BitSlice2_out1                   : std_logic;
  SIGNAL BitSlice4_out1_1                 : std_logic;
  SIGNAL C4_out1                          : unsigned(7 DOWNTO 0);
  SIGNAL Sum_0_out1                       : std_logic;
  SIGNAL exp_a_cor_shift_length_out1      : unsigned(7 DOWNTO 0);
  SIGNAL C2_out1                          : unsigned(7 DOWNTO 0);
  SIGNAL if_shift_length_exp_a_cor_out1   : unsigned(7 DOWNTO 0);
  SIGNAL BitSlice2_out1_1                 : std_logic;
  SIGNAL C3_out1                          : unsigned(7 DOWNTO 0);
  SIGNAL if_Sum_0_out1                    : unsigned(7 DOWNTO 0);
  SIGNAL if_bitget_Sum_Sum_WordLength_1_out1 : unsigned(7 DOWNTO 0);
  SIGNAL C_out1_2                         : unsigned(7 DOWNTO 0);
  SIGNAL exp_a_cor_1_out1_1               : unsigned(7 DOWNTO 0);
  SIGNAL if_bitget_Sum_Sum_WordLength_1_out1_1 : unsigned(7 DOWNTO 0);
  SIGNAL Delay14_out1                     : unsigned(7 DOWNTO 0);
  SIGNAL if_bitget_Sum_Sum_WordLength_out1_1 : unsigned(7 DOWNTO 0);
  SIGNAL cast_1_like_Exp_out1             : unsigned(7 DOWNTO 0);
  SIGNAL Exp_cast_1_like_Exp_out1         : unsigned(7 DOWNTO 0);
  SIGNAL if_bitget_Mant_tmp_Mant_tmp_Wor_out1 : unsigned(7 DOWNTO 0);
  SIGNAL Exponent_0_out1_2                : std_logic;
  SIGNAL BitSlice3_out1_1                 : unsigned(22 DOWNTO 0);
  SIGNAL Mantissa_0_out1                  : std_logic;
  SIGNAL alphaExponent_0_Mantissa_out1    : std_logic;
  SIGNAL Constant_out1_2                  : std_logic;
  SIGNAL Switch_out1_1                    : std_logic;
  SIGNAL Delay12_out1_1                   : std_logic;
  SIGNAL Delay29_out1                     : std_logic;
  SIGNAL Delay14_reg_rsvd                 : std_logic_vector(0 TO 1);
  SIGNAL Delay14_reg_next                 : std_logic_vector(0 TO 1);
  SIGNAL Delay14_out1_1                   : std_logic;
  SIGNAL alphaaSign_1_bSign_1_out1        : std_logic;
  SIGNAL Delay9_out1                      : std_logic;
  SIGNAL Delay25_out1                     : std_logic;
  SIGNAL Delay13_reg_rsvd                 : std_logic_vector(0 TO 1);
  SIGNAL Delay13_reg_next                 : std_logic_vector(0 TO 1);
  SIGNAL Delay13_out1_1                   : std_logic;
  SIGNAL if_Exponent_0_Mantissa_out1      : std_logic;
  SIGNAL Delay6_out1                      : std_logic;
  SIGNAL Delay32_out1                     : unsigned(7 DOWNTO 0);
  SIGNAL Delay34_out1                     : unsigned(7 DOWNTO 0);
  SIGNAL Delay15_reg_rsvd                 : vector_of_unsigned8(0 TO 1);
  SIGNAL Delay15_reg_next                 : vector_of_unsigned8(0 TO 1);
  SIGNAL Delay15_out1_1                   : unsigned(7 DOWNTO 0);
  SIGNAL if_aExponent_cfType_Exponent_out1 : unsigned(7 DOWNTO 0);
  SIGNAL Delay7_out1                      : unsigned(7 DOWNTO 0);
  SIGNAL opp_signs_exp_b_cfType_out1      : std_logic;
  SIGNAL mant_a_0_out1                    : std_logic;
  SIGNAL alphamant_a_0_opp_signs_out1     : std_logic;
  SIGNAL BitSet_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL if_mant_a_0_opp_signs_out1       : unsigned(22 DOWNTO 0);
  SIGNAL Delay2_out1_3                    : unsigned(22 DOWNTO 0);
  SIGNAL Delay38_out1                     : unsigned(22 DOWNTO 0);
  SIGNAL Delay17_reg_rsvd                 : vector_of_unsigned23(0 TO 1);
  SIGNAL Delay17_reg_next                 : vector_of_unsigned23(0 TO 1);
  SIGNAL Delay17_out1                     : unsigned(22 DOWNTO 0);
  SIGNAL if_aExponent_cfType_Exponent_1_out1 : unsigned(22 DOWNTO 0);
  SIGNAL Delay8_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL nfp_out_pack                     : unsigned(31 DOWNTO 0);

BEGIN
  nfp_in1_unsigned <= unsigned(nfp_in1);

  -- Split 32 bit word into FP sign, exponent, mantissa
  AS <= nfp_in1_unsigned(31);
  AE <= nfp_in1_unsigned(30 DOWNTO 23);
  AM <= nfp_in1_unsigned(22 DOWNTO 0);

  Delay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay1_out1 <= AE;
      END IF;
    END IF;
  END PROCESS Delay1_process;


  nfp_in2_unsigned <= unsigned(nfp_in2);

  -- Split 32 bit word into FP sign, exponent, mantissa
  BS <= nfp_in2_unsigned(31);
  BE <= nfp_in2_unsigned(30 DOWNTO 23);
  BM <= nfp_in2_unsigned(22 DOWNTO 0);

  Delay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay4_out1 <= BE;
      END IF;
    END IF;
  END PROCESS Delay4_process;


  
  Relational_Operator1_relop1 <= '1' WHEN Delay1_out1 = Delay4_out1 ELSE
      '0';

  Delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay2_out1 <= AM;
      END IF;
    END IF;
  END PROCESS Delay2_process;


  Delay5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay5_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay5_out1 <= BM;
      END IF;
    END IF;
  END PROCESS Delay5_process;


  
  Relational_Operator_relop1 <= '1' WHEN Delay1_out1 > Delay4_out1 ELSE
      '0';

  
  bitconcat_aExponent_aMantissa_relop1 <= '1' WHEN Delay2_out1 >= Delay5_out1 ELSE
      '0';

  Logical_Operator_out1 <= Relational_Operator1_relop1 AND bitconcat_aExponent_aMantissa_relop1;

  Logical_Operator1_out1 <= Relational_Operator_relop1 OR Logical_Operator_out1;

  
  if_bitconcat_aExponent_aMantiss_out1 <= Delay4_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay1_out1;

  
  aExponent_cfType_Exponent_I_out1 <= '1' WHEN if_bitconcat_aExponent_aMantiss_out1 = to_unsigned(16#FF#, 8) 
    ELSE
      '0';

  Delay11_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay11_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay11_out1 <= aExponent_cfType_Exponent_I_out1;
      END IF;
    END IF;
  END PROCESS Delay11_process;


  Delay42_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay42_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay42_out1 <= Delay11_out1;
      END IF;
    END IF;
  END PROCESS Delay42_process;


  Delay18_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay18_reg_rsvd(0) <= '0';
        Delay18_reg_rsvd(1) <= '0';
      ELSIF enb = '1' THEN
        Delay18_reg_rsvd(0) <= Delay18_reg_next(0);
        Delay18_reg_rsvd(1) <= Delay18_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay18_process;

  Delay18_out1 <= Delay18_reg_rsvd(1);
  Delay18_reg_next(0) <= Delay42_out1;
  Delay18_reg_next(1) <= Delay18_reg_rsvd(0);

  
  Exponent_0_out1 <= '1' WHEN if_bitconcat_aExponent_aMantiss_out1 = to_unsigned(16#00#, 8) ELSE
      '0';

  C_out1 <= to_unsigned(16#01#, 8);

  
  if_Exponent_0_out1 <= if_bitconcat_aExponent_aMantiss_out1 WHEN Exponent_0_out1 = '0' ELSE
      C_out1;

  Delay_rsvd_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay_out1 <= if_Exponent_0_out1;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_process;


  Delay4_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay4_out1_1 <= Delay_out1;
      END IF;
    END IF;
  END PROCESS Delay4_1_process;


  Delay2_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay2_out1_1 <= Delay4_out1_1;
      END IF;
    END IF;
  END PROCESS Delay2_1_process;


  
  exp_norm_cfType_Exponent_In_out1 <= '1' WHEN Delay2_out1_1 = to_unsigned(16#FE#, 8) ELSE
      '0';

  alphaExponent_0_cfType_Exp_out1 <= aExponent_cfType_Exponent_I_out1 OR Exponent_0_out1;

  alpha1_out1 <= to_unsigned(16#1#, 3);

  alpha0_out1 <= to_unsigned(16#0#, 3);

  
  if_Exponent_0_cfType_Exp_out1 <= alpha1_out1 WHEN alphaExponent_0_cfType_Exp_out1 = '0' ELSE
      alpha0_out1;

  
  if_bitconcat_aExponent_aMantiss_1_ou_1 <= Delay5_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay2_out1;

  Bit_Concat_out1 <= if_Exponent_0_cfType_Exp_out1 & if_bitconcat_aExponent_aMantiss_1_ou_1;

  alpha0_1_out1 <= to_unsigned(16#0#, 2);

  Bit_Concat1_out1 <= Bit_Concat_out1 & alpha0_1_out1;

  Data_Type_Conversion_out1 <= signed(Bit_Concat1_out1);

  Delay2_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_2 <= to_signed(16#0000000#, 28);
      ELSIF enb = '1' THEN
        Delay2_out1_2 <= Data_Type_Conversion_out1;
      END IF;
    END IF;
  END PROCESS Delay2_2_process;


  Delay5_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay5_out1_1 <= to_signed(16#0000000#, 28);
      ELSIF enb = '1' THEN
        Delay5_out1_1 <= Delay2_out1_2;
      END IF;
    END IF;
  END PROCESS Delay5_1_process;


  Delay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay3_out1 <= BS;
      END IF;
    END IF;
  END PROCESS Delay3_process;


  Logical_Operator_out1_1 <=  NOT Delay3_out1;

  Delay_rsvd_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1_1 <= '0';
      ELSIF enb = '1' THEN
        Delay_out1_1 <= AS;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_1_process;


  
  if_bitconcat_aExponent_aMantiss_2_ou_1 <= Logical_Operator_out1_1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay_out1_1;

  
  if_bitconcat_aExponent_aMantiss_5_ou_1 <= Delay_out1_1 WHEN Logical_Operator1_out1 = '0' ELSE
      Logical_Operator_out1_1;

  bitxor_out1 <= if_bitconcat_aExponent_aMantiss_2_ou_1 XOR if_bitconcat_aExponent_aMantiss_5_ou_1;

  Delay10_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay10_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay10_out1 <= bitxor_out1;
      END IF;
    END IF;
  END PROCESS Delay10_process;


  
  if_bitconcat_aExponent_aMantiss_3_ou_1 <= Delay1_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay4_out1;

  
  exp_b_cfType_Exponent_Inf_o_out1 <= '1' WHEN if_bitconcat_aExponent_aMantiss_3_ou_1 = to_unsigned(16#FF#, 
    8) ELSE
      '0';

  
  Exponent_0_out1_1 <= '1' WHEN if_bitconcat_aExponent_aMantiss_3_ou_1 = to_unsigned(16#00#, 8) ELSE
      '0';

  alphaExponent_0_cfType_Exp_out1_1 <= exp_b_cfType_Exponent_Inf_o_out1 OR Exponent_0_out1_1;

  alpha1_out1_1 <= to_unsigned(16#1#, 3);

  alpha0_out1_1 <= to_unsigned(16#0#, 3);

  
  if_Exponent_0_cfType_Exp_out1_1 <= alpha1_out1_1 WHEN alphaExponent_0_cfType_Exp_out1_1 = '0' ELSE
      alpha0_out1_1;

  
  if_bitconcat_aExponent_aMantiss_4_ou_1 <= Delay2_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay5_out1;

  Bit_Concat_out1_1 <= if_Exponent_0_cfType_Exp_out1_1 & if_bitconcat_aExponent_aMantiss_4_ou_1;

  alpha0_1_out1_1 <= to_unsigned(16#0#, 2);

  Bit_Concat1_out1_1 <= Bit_Concat_out1_1 & alpha0_1_out1_1;

  Data_Type_Conversion_out1_1 <= signed(Bit_Concat1_out1_1);

  Delay1_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_1 <= to_signed(16#0000000#, 28);
      ELSIF enb = '1' THEN
        Delay1_out1_1 <= Data_Type_Conversion_out1_1;
      END IF;
    END IF;
  END PROCESS Delay1_1_process;


  alphamant_b_ext_in0 <=  - (resize(Delay1_out1_1, 29));
  alphamant_b_ext_out1 <= alphamant_b_ext_in0(27 DOWNTO 0);

  
  if_opp_Sign_out1 <= Delay1_out1_1 WHEN Delay10_out1 = '0' ELSE
      alphamant_b_ext_out1;

  C_out1_1 <= to_unsigned(16#01#, 8);

  
  if_Exponent_0_out1_1 <= if_bitconcat_aExponent_aMantiss_3_ou_1 WHEN Exponent_0_out1_1 = '0' ELSE
      C_out1_1;

  Delay_rsvd_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1_2 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay_out1_2 <= if_Exponent_0_out1_1;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_2_process;


  storedInteger_exp_a_cor_sto_sub_cast <= signed(resize(Delay_out1, 32));
  storedInteger_exp_a_cor_sto_sub_cast_1 <= signed(resize(Delay_out1_2, 32));
  storedInteger_exp_a_cor_sto_out1 <= storedInteger_exp_a_cor_sto_sub_cast - 
    storedInteger_exp_a_cor_sto_sub_cast_1;

  Bit_Slice2_out1 <= unsigned(storedInteger_exp_a_cor_sto_out1(7 DOWNTO 5));

  
  Compare_To_Zero_out1 <= '1' WHEN Bit_Slice2_out1 = to_unsigned(16#0#, 3) ELSE
      '0';

  Constant_out1 <= to_unsigned(16#1F#, 5);

  Bit_Slice_out1 <= unsigned(storedInteger_exp_a_cor_sto_out1(4 DOWNTO 0));

  
  if_opp_Sign_1_out1 <= Constant_out1 WHEN Compare_To_Zero_out1 = '0' ELSE
      Bit_Slice_out1;

  bitsra_mant_b_ext_shift_lengt_out1 <= SHIFT_RIGHT(if_opp_Sign_out1, to_integer(if_opp_Sign_1_out1));

  Delay1_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_2 <= to_signed(16#0000000#, 28);
      ELSIF enb = '1' THEN
        Delay1_out1_2 <= bitsra_mant_b_ext_shift_lengt_out1;
      END IF;
    END IF;
  END PROCESS Delay1_2_process;


  mant_a_ext_mant_b_shifted_add_temp <= resize(Delay5_out1_1, 32) + resize(Delay1_out1_2, 32);
  mant_a_ext_mant_b_shifted_out1 <= unsigned(mant_a_ext_mant_b_shifted_add_temp(26 DOWNTO 0));

  BitSlice_out1 <= mant_a_ext_mant_b_shifted_out1(26);

  Delay3_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1_1 <= '0';
      ELSIF enb = '1' THEN
        Delay3_out1_1 <= BitSlice_out1;
      END IF;
    END IF;
  END PROCESS Delay3_1_process;


  Logical_Operator_out1_2 <= exp_norm_cfType_Exponent_In_out1 AND Delay3_out1_1;

  Delay13_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay13_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay13_out1 <= Logical_Operator_out1_2;
      END IF;
    END IF;
  END PROCESS Delay13_process;


  Delay1_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_3 <= to_unsigned(16#0000000#, 27);
      ELSIF enb = '1' THEN
        Delay1_out1_3 <= mant_a_ext_mant_b_shifted_out1;
      END IF;
    END IF;
  END PROCESS Delay1_3_process;


  BitSlice3_out1 <= mant_a_ext_mant_b_shifted_out1(25 DOWNTO 0);

  Bit_Slice5_out1 <= BitSlice3_out1(25);

  Bit_Slice3_out1 <= BitSlice3_out1(24);

  Logical_Operator1_out1_1 <= Bit_Slice5_out1 OR Bit_Slice3_out1;

  Bit_Slice2_out1_1 <= BitSlice3_out1(23 DOWNTO 16);

  Bit_Slice16_out1 <= Bit_Slice2_out1_1(7);

  Bit_Slice15_out1 <= Bit_Slice2_out1_1(6);

  Logical_Operator5_out1 <= Bit_Slice16_out1 OR Bit_Slice15_out1;

  Bit_Slice14_out1 <= Bit_Slice2_out1_1(5);

  Bit_Slice13_out1 <= Bit_Slice2_out1_1(4);

  Logical_Operator7_out1 <= Bit_Slice14_out1 OR Bit_Slice13_out1;

  Logical_Operator6_out1 <= Logical_Operator5_out1 OR Logical_Operator7_out1;

  Bit_Slice12_out1 <= Bit_Slice2_out1_1(3);

  Bit_Slice11_out1 <= Bit_Slice2_out1_1(2);

  Logical_Operator4_out1 <= Bit_Slice12_out1 OR Bit_Slice11_out1;

  Bit_Slice10_out1 <= Bit_Slice2_out1_1(1);

  Bit_Slice9_out1 <= Bit_Slice2_out1_1(0);

  Logical_Operator14_out1 <= Bit_Slice10_out1 OR Bit_Slice9_out1;

  Logical_Operator13_out1 <= Logical_Operator4_out1 OR Logical_Operator14_out1;

  Logical_Operator12_out1 <= Logical_Operator6_out1 OR Logical_Operator13_out1;

  Bit_Slice1_out1 <= BitSlice3_out1(15 DOWNTO 8);

  Bit_Slice16_out1_1 <= Bit_Slice1_out1(7);

  Bit_Slice15_out1_1 <= Bit_Slice1_out1(6);

  Logical_Operator5_out1_1 <= Bit_Slice16_out1_1 OR Bit_Slice15_out1_1;

  Bit_Slice14_out1_1 <= Bit_Slice1_out1(5);

  Bit_Slice13_out1_1 <= Bit_Slice1_out1(4);

  Logical_Operator7_out1_1 <= Bit_Slice14_out1_1 OR Bit_Slice13_out1_1;

  Logical_Operator6_out1_1 <= Logical_Operator5_out1_1 OR Logical_Operator7_out1_1;

  Bit_Slice12_out1_1 <= Bit_Slice1_out1(3);

  Bit_Slice11_out1_1 <= Bit_Slice1_out1(2);

  Logical_Operator4_out1_1 <= Bit_Slice12_out1_1 OR Bit_Slice11_out1_1;

  Bit_Slice10_out1_1 <= Bit_Slice1_out1(1);

  Bit_Slice9_out1_1 <= Bit_Slice1_out1(0);

  Logical_Operator14_out1_1 <= Bit_Slice10_out1_1 OR Bit_Slice9_out1_1;

  Logical_Operator13_out1_1 <= Logical_Operator4_out1_1 OR Logical_Operator14_out1_1;

  Bit_Slice4_out1 <= BitSlice3_out1(7 DOWNTO 0);

  Bit_Slice8_out1 <= Bit_Slice4_out1(7);

  Bit_Slice7_out1 <= Bit_Slice4_out1(6);

  Logical_Operator1_out1_2 <= Bit_Slice8_out1 OR Bit_Slice7_out1;

  Bit_Slice6_out1 <= Bit_Slice4_out1(5);

  Bit_Slice5_out1_1 <= Bit_Slice4_out1(4);

  Logical_Operator3_out1 <= Bit_Slice6_out1 OR Bit_Slice5_out1_1;

  Bit_Slice3_out1_1 <= Bit_Slice4_out1(3);

  Bit_Slice2_out1_2 <= Bit_Slice4_out1(2);

  Bit_Slice1_out1_1 <= Bit_Slice4_out1(1);

  Bit_Slice_out1_1 <= Bit_Slice4_out1(0);

  Constant_out1_1 <= to_unsigned(16#1A#, 5);

  Constant1_out1 <= to_unsigned(16#19#, 5);

  
  Switch_out1 <= Constant_out1_1 WHEN Bit_Slice_out1_1 = '0' ELSE
      Constant1_out1;

  Logical_Operator_out1_3 <= Bit_Slice3_out1_1 OR Bit_Slice2_out1_2;

  Constant2_out1 <= to_unsigned(16#18#, 5);

  
  Switch1_out1 <= Switch_out1 WHEN Bit_Slice1_out1_1 = '0' ELSE
      Constant2_out1;

  Constant3_out1 <= to_unsigned(16#17#, 5);

  
  Switch2_out1 <= Constant_out1_1 WHEN Bit_Slice2_out1_2 = '0' ELSE
      Constant3_out1;

  Constant4_out1 <= to_unsigned(16#16#, 5);

  Logical_Operator2_out1 <= Logical_Operator1_out1_2 OR Logical_Operator3_out1;

  
  Switch3_out1 <= Switch2_out1 WHEN Bit_Slice3_out1_1 = '0' ELSE
      Constant4_out1;

  
  Switch4_out1 <= Switch1_out1 WHEN Logical_Operator_out1_3 = '0' ELSE
      Switch3_out1;

  Constant5_out1 <= to_unsigned(16#15#, 5);

  
  Switch5_out1 <= Constant_out1_1 WHEN Bit_Slice5_out1_1 = '0' ELSE
      Constant5_out1;

  Constant6_out1 <= to_unsigned(16#14#, 5);

  
  Switch6_out1 <= Switch5_out1 WHEN Bit_Slice6_out1 = '0' ELSE
      Constant6_out1;

  Constant7_out1 <= to_unsigned(16#13#, 5);

  
  Switch7_out1 <= Constant_out1_1 WHEN Bit_Slice7_out1 = '0' ELSE
      Constant7_out1;

  Constant8_out1 <= to_unsigned(16#12#, 5);

  
  Switch8_out1 <= Switch7_out1 WHEN Bit_Slice8_out1 = '0' ELSE
      Constant8_out1;

  Logical_Operator12_out1_1 <= Logical_Operator6_out1_1 OR Logical_Operator13_out1_1;

  
  Switch9_out1 <= Switch6_out1 WHEN Logical_Operator1_out1_2 = '0' ELSE
      Switch8_out1;

  
  Switch10_out1 <= Switch4_out1 WHEN Logical_Operator2_out1 = '0' ELSE
      Switch9_out1;

  Constant9_out1 <= to_unsigned(16#11#, 5);

  
  Switch11_out1 <= Constant_out1_1 WHEN Bit_Slice9_out1_1 = '0' ELSE
      Constant9_out1;

  Constant10_out1 <= to_unsigned(16#10#, 5);

  
  Switch12_out1 <= Switch11_out1 WHEN Bit_Slice10_out1_1 = '0' ELSE
      Constant10_out1;

  Constant11_out1 <= to_unsigned(16#0F#, 5);

  
  Switch14_out1 <= Constant_out1_1 WHEN Bit_Slice11_out1_1 = '0' ELSE
      Constant11_out1;

  Constant12_out1 <= to_unsigned(16#0E#, 5);

  
  Switch15_out1 <= Switch14_out1 WHEN Bit_Slice12_out1_1 = '0' ELSE
      Constant12_out1;

  
  Switch16_out1 <= Switch12_out1 WHEN Logical_Operator4_out1_1 = '0' ELSE
      Switch15_out1;

  Constant13_out1 <= to_unsigned(16#0D#, 5);

  
  Switch17_out1 <= Constant_out1_1 WHEN Bit_Slice13_out1_1 = '0' ELSE
      Constant13_out1;

  Constant14_out1 <= to_unsigned(16#0C#, 5);

  
  Switch18_out1 <= Switch17_out1 WHEN Bit_Slice14_out1_1 = '0' ELSE
      Constant14_out1;

  Constant15_out1 <= to_unsigned(16#0B#, 5);

  
  Switch19_out1 <= Constant_out1_1 WHEN Bit_Slice15_out1_1 = '0' ELSE
      Constant15_out1;

  Constant16_out1 <= to_unsigned(16#0A#, 5);

  
  Switch20_out1 <= Switch19_out1 WHEN Bit_Slice16_out1_1 = '0' ELSE
      Constant16_out1;

  
  Switch21_out1 <= Switch18_out1 WHEN Logical_Operator5_out1_1 = '0' ELSE
      Switch20_out1;

  Logical_Operator_out1_4 <= Logical_Operator1_out1_1 OR Logical_Operator12_out1;

  
  Switch13_out1 <= Switch16_out1 WHEN Logical_Operator6_out1_1 = '0' ELSE
      Switch21_out1;

  
  Switch33_out1 <= Switch10_out1 WHEN Logical_Operator12_out1_1 = '0' ELSE
      Switch13_out1;

  Constant9_out1_1 <= to_unsigned(16#09#, 5);

  
  Switch11_out1_1 <= Constant_out1_1 WHEN Bit_Slice9_out1 = '0' ELSE
      Constant9_out1_1;

  Constant10_out1_1 <= to_unsigned(16#08#, 5);

  
  Switch12_out1_1 <= Switch11_out1_1 WHEN Bit_Slice10_out1 = '0' ELSE
      Constant10_out1_1;

  Constant11_out1_1 <= to_unsigned(16#07#, 5);

  
  Switch14_out1_1 <= Constant_out1_1 WHEN Bit_Slice11_out1 = '0' ELSE
      Constant11_out1_1;

  Constant12_out1_1 <= to_unsigned(16#06#, 5);

  
  Switch15_out1_1 <= Switch14_out1_1 WHEN Bit_Slice12_out1 = '0' ELSE
      Constant12_out1_1;

  
  Switch16_out1_1 <= Switch12_out1_1 WHEN Logical_Operator4_out1 = '0' ELSE
      Switch15_out1_1;

  Constant13_out1_1 <= to_unsigned(16#05#, 5);

  
  Switch17_out1_1 <= Constant_out1_1 WHEN Bit_Slice13_out1 = '0' ELSE
      Constant13_out1_1;

  Constant14_out1_1 <= to_unsigned(16#04#, 5);

  
  Switch18_out1_1 <= Switch17_out1_1 WHEN Bit_Slice14_out1 = '0' ELSE
      Constant14_out1_1;

  Constant15_out1_1 <= to_unsigned(16#03#, 5);

  
  Switch19_out1_1 <= Constant_out1_1 WHEN Bit_Slice15_out1 = '0' ELSE
      Constant15_out1_1;

  Constant16_out1_1 <= to_unsigned(16#02#, 5);

  
  Switch20_out1_1 <= Switch19_out1_1 WHEN Bit_Slice16_out1 = '0' ELSE
      Constant16_out1_1;

  
  Switch21_out1_1 <= Switch18_out1_1 WHEN Logical_Operator5_out1 = '0' ELSE
      Switch20_out1_1;

  
  Switch13_out1_1 <= Switch16_out1_1 WHEN Logical_Operator6_out1 = '0' ELSE
      Switch21_out1_1;

  Constant1_out1_1 <= to_unsigned(16#01#, 5);

  
  Switch3_out1_1 <= Constant_out1_1 WHEN Bit_Slice3_out1 = '0' ELSE
      Constant1_out1_1;

  Constant2_out1_1 <= to_unsigned(16#00#, 5);

  
  Switch2_out1_1 <= Switch3_out1_1 WHEN Bit_Slice5_out1 = '0' ELSE
      Constant2_out1_1;

  
  Switch1_out1_1 <= Switch13_out1_1 WHEN Logical_Operator1_out1_1 = '0' ELSE
      Switch2_out1_1;

  
  Switch34_out1 <= Switch33_out1 WHEN Logical_Operator_out1_4 = '0' ELSE
      Switch1_out1_1;

  Delay_rsvd_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1_3 <= to_unsigned(16#00#, 5);
      ELSIF enb = '1' THEN
        Delay_out1_3 <= Switch34_out1;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_3_process;


  Bit_Slice_out1_2 <= Delay2_out1_1(4 DOWNTO 0);

  
  shift_length_exp_a_cor_relop1 <= '1' WHEN Delay_out1_3 >= Bit_Slice_out1_2 ELSE
      '0';

  Bit_Slice1_out1_2 <= Delay2_out1_1(7 DOWNTO 5);

  
  Compare_To_Zero_out1_1 <= '1' WHEN Bit_Slice1_out1_2 = to_unsigned(16#0#, 3) ELSE
      '0';

  Logical_Operator1_out1_3 <= shift_length_exp_a_cor_relop1 AND Compare_To_Zero_out1_1;

  C1_out1 <= to_unsigned(16#01#, 8);

  exp_a_cor_1_out1 <= Bit_Slice_out1_2 - resize(C1_out1, 5);

  
  if_shift_length_exp_a_cor_1_out1 <= Delay_out1_3 WHEN Logical_Operator1_out1_3 = '0' ELSE
      exp_a_cor_1_out1;

  bitsll_Sum_shift_length_out1 <= Delay1_out1_3 sll to_integer(if_shift_length_exp_a_cor_1_out1);

  bitsrl_Sum_1_out1 <= Delay1_out1_3 srl 1;

  
  if_bitget_Sum_Sum_WordLength_out1 <= bitsll_Sum_shift_length_out1 WHEN Delay3_out1_1 = '0' ELSE
      bitsrl_Sum_1_out1;

  Delay15_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay15_out1 <= to_unsigned(16#0000000#, 27);
      ELSIF enb = '1' THEN
        Delay15_out1 <= if_bitget_Sum_Sum_WordLength_out1;
      END IF;
    END IF;
  END PROCESS Delay15_process;


  C5_out1 <= to_unsigned(16#0000000#, 27);

  
  if_exp_norm_cfType_Exponent_I_out1 <= Delay15_out1 WHEN Delay13_out1 = '0' ELSE
      C5_out1;

  BitSlice6_out1 <= if_exp_norm_cfType_Exponent_I_out1(24 DOWNTO 1);

  BitSlice5_out1 <= if_exp_norm_cfType_Exponent_I_out1(0);

  Bit_Slice13_out1_2 <= if_opp_Sign_1_out1(4);

  Bit_Slice12_out1_2 <= if_opp_Sign_1_out1(3);

  Bit_Slice10_out1_2 <= if_opp_Sign_1_out1(2);

  Bit_Slice11_out1_2 <= if_opp_Sign_1_out1(1);

  Bit_Slice14_out1_2 <= if_opp_Sign_1_out1(0);

  Bit_Slice7_out1_1 <= unsigned(if_opp_Sign_out1(2 DOWNTO 0));

  Constant1_out1_2 <= '0';

  Bit_Concat_out1_2 <= Bit_Slice7_out1_1 & Constant1_out1_2;

  Bit_Slice_out1_3 <= Bit_Concat_out1_2(0);

  Data_Type_Conversion_out1_2 <= Bit_Slice_out1_3;

  Bit_Slice1_out1_3 <= Bit_Concat_out1_2(1);

  Logical_Operator_out1_5 <= Bit_Slice1_out1_3 OR Data_Type_Conversion_out1_2;

  
  Switch6_out1_1 <= Data_Type_Conversion_out1_2 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_5;

  Bit_Slice2_out1_3 <= Bit_Concat_out1_2(2);

  Logical_Operator1_out1_4 <= Bit_Slice2_out1_3 OR Logical_Operator_out1_5;

  Bit_Slice3_out1_2 <= Bit_Concat_out1_2(3);

  Logical_Operator2_out1_1 <= Bit_Slice3_out1_2 OR Logical_Operator1_out1_4;

  
  Switch7_out1_1 <= Logical_Operator1_out1_4 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_1;

  
  Switch3_out1_2 <= Switch6_out1_1 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_1;

  Bit_Slice8_out1_1 <= unsigned(if_opp_Sign_out1(6 DOWNTO 3));

  Bit_Slice_out1_4 <= Bit_Slice8_out1_1(0);

  Logical_Operator3_out1_1 <= Bit_Slice_out1_4 OR Logical_Operator2_out1_1;

  Bit_Slice1_out1_4 <= Bit_Slice8_out1_1(1);

  Logical_Operator_out1_6 <= Bit_Slice1_out1_4 OR Logical_Operator3_out1_1;

  
  Switch6_out1_2 <= Logical_Operator3_out1_1 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_6;

  Bit_Slice2_out1_4 <= Bit_Slice8_out1_1(2);

  Logical_Operator1_out1_5 <= Bit_Slice2_out1_4 OR Logical_Operator_out1_6;

  Bit_Slice3_out1_3 <= Bit_Slice8_out1_1(3);

  Logical_Operator2_out1_2 <= Bit_Slice3_out1_3 OR Logical_Operator1_out1_5;

  
  Switch7_out1_2 <= Logical_Operator1_out1_5 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_2;

  
  Switch3_out1_3 <= Switch6_out1_2 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_2;

  
  Switch6_out1_3 <= Switch3_out1_2 WHEN Bit_Slice10_out1_2 = '0' ELSE
      Switch3_out1_3;

  Bit_Slice9_out1_2 <= unsigned(if_opp_Sign_out1(10 DOWNTO 7));

  Bit_Slice_out1_5 <= Bit_Slice9_out1_2(0);

  Logical_Operator3_out1_2 <= Bit_Slice_out1_5 OR Logical_Operator2_out1_2;

  Bit_Slice1_out1_5 <= Bit_Slice9_out1_2(1);

  Logical_Operator_out1_7 <= Bit_Slice1_out1_5 OR Logical_Operator3_out1_2;

  
  Switch6_out1_4 <= Logical_Operator3_out1_2 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_7;

  Bit_Slice2_out1_5 <= Bit_Slice9_out1_2(2);

  Logical_Operator1_out1_6 <= Bit_Slice2_out1_5 OR Logical_Operator_out1_7;

  Bit_Slice3_out1_4 <= Bit_Slice9_out1_2(3);

  Logical_Operator2_out1_3 <= Bit_Slice3_out1_4 OR Logical_Operator1_out1_6;

  
  Switch7_out1_3 <= Logical_Operator1_out1_6 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_3;

  
  Switch3_out1_4 <= Switch6_out1_4 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_3;

  Bit_Slice3_out1_5 <= unsigned(if_opp_Sign_out1(14 DOWNTO 11));

  Bit_Slice_out1_6 <= Bit_Slice3_out1_5(0);

  Logical_Operator3_out1_3 <= Bit_Slice_out1_6 OR Logical_Operator2_out1_3;

  Bit_Slice1_out1_6 <= Bit_Slice3_out1_5(1);

  Logical_Operator_out1_8 <= Bit_Slice1_out1_6 OR Logical_Operator3_out1_3;

  
  Switch6_out1_5 <= Logical_Operator3_out1_3 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_8;

  Bit_Slice2_out1_6 <= Bit_Slice3_out1_5(2);

  Logical_Operator1_out1_7 <= Bit_Slice2_out1_6 OR Logical_Operator_out1_8;

  Bit_Slice3_out1_6 <= Bit_Slice3_out1_5(3);

  Logical_Operator2_out1_4 <= Bit_Slice3_out1_6 OR Logical_Operator1_out1_7;

  
  Switch7_out1_4 <= Logical_Operator1_out1_7 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_4;

  
  Switch3_out1_5 <= Switch6_out1_5 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_4;

  
  Switch7_out1_5 <= Switch3_out1_4 WHEN Bit_Slice10_out1_2 = '0' ELSE
      Switch3_out1_5;

  
  Switch3_out1_6 <= Switch6_out1_3 WHEN Bit_Slice12_out1_2 = '0' ELSE
      Switch7_out1_5;

  Bit_Slice4_out1_1 <= unsigned(if_opp_Sign_out1(18 DOWNTO 15));

  Bit_Slice_out1_7 <= Bit_Slice4_out1_1(0);

  Logical_Operator3_out1_4 <= Bit_Slice_out1_7 OR Logical_Operator2_out1_4;

  Bit_Slice1_out1_7 <= Bit_Slice4_out1_1(1);

  Logical_Operator_out1_9 <= Bit_Slice1_out1_7 OR Logical_Operator3_out1_4;

  
  Switch6_out1_6 <= Logical_Operator3_out1_4 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_9;

  Bit_Slice2_out1_7 <= Bit_Slice4_out1_1(2);

  Logical_Operator1_out1_8 <= Bit_Slice2_out1_7 OR Logical_Operator_out1_9;

  Bit_Slice3_out1_7 <= Bit_Slice4_out1_1(3);

  Logical_Operator2_out1_5 <= Bit_Slice3_out1_7 OR Logical_Operator1_out1_8;

  
  Switch7_out1_6 <= Logical_Operator1_out1_8 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_5;

  
  Switch3_out1_7 <= Switch6_out1_6 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_6;

  Bit_Slice5_out1_2 <= unsigned(if_opp_Sign_out1(22 DOWNTO 19));

  Bit_Slice_out1_8 <= Bit_Slice5_out1_2(0);

  Logical_Operator3_out1_5 <= Bit_Slice_out1_8 OR Logical_Operator2_out1_5;

  Bit_Slice1_out1_8 <= Bit_Slice5_out1_2(1);

  Logical_Operator_out1_10 <= Bit_Slice1_out1_8 OR Logical_Operator3_out1_5;

  
  Switch6_out1_7 <= Logical_Operator3_out1_5 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_10;

  Bit_Slice2_out1_8 <= Bit_Slice5_out1_2(2);

  Logical_Operator1_out1_9 <= Bit_Slice2_out1_8 OR Logical_Operator_out1_10;

  Bit_Slice3_out1_8 <= Bit_Slice5_out1_2(3);

  Logical_Operator2_out1_6 <= Bit_Slice3_out1_8 OR Logical_Operator1_out1_9;

  
  Switch7_out1_7 <= Logical_Operator1_out1_9 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_6;

  
  Switch3_out1_8 <= Switch6_out1_7 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_7;

  
  Switch6_out1_8 <= Switch3_out1_7 WHEN Bit_Slice10_out1_2 = '0' ELSE
      Switch3_out1_8;

  Bit_Slice6_out1_1 <= unsigned(if_opp_Sign_out1(26 DOWNTO 23));

  Bit_Slice_out1_9 <= Bit_Slice6_out1_1(0);

  Logical_Operator3_out1_6 <= Bit_Slice_out1_9 OR Logical_Operator2_out1_6;

  Bit_Slice1_out1_9 <= Bit_Slice6_out1_1(1);

  Logical_Operator_out1_11 <= Bit_Slice1_out1_9 OR Logical_Operator3_out1_6;

  
  Switch6_out1_9 <= Logical_Operator3_out1_6 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator_out1_11;

  Bit_Slice2_out1_9 <= Bit_Slice6_out1_1(2);

  Logical_Operator1_out1_10 <= Bit_Slice2_out1_9 OR Logical_Operator_out1_11;

  Bit_Slice3_out1_9 <= Bit_Slice6_out1_1(3);

  Logical_Operator2_out1_7 <= Bit_Slice3_out1_9 OR Logical_Operator1_out1_10;

  
  Switch7_out1_8 <= Logical_Operator1_out1_10 WHEN Bit_Slice14_out1_2 = '0' ELSE
      Logical_Operator2_out1_7;

  
  Switch3_out1_9 <= Switch6_out1_9 WHEN Bit_Slice11_out1_2 = '0' ELSE
      Switch7_out1_8;

  Bit_Slice1_out1_10 <= if_opp_Sign_out1(27);

  Logical_Operator_out1_12 <=  NOT Bit_Slice1_out1_10;

  Logical_Operator1_out1_11 <= Logical_Operator_out1_12 AND Logical_Operator2_out1_7;

  
  Switch7_out1_9 <= Switch3_out1_9 WHEN Bit_Slice10_out1_2 = '0' ELSE
      Logical_Operator1_out1_11;

  
  Switch3_out1_10 <= Switch6_out1_8 WHEN Bit_Slice12_out1_2 = '0' ELSE
      Switch7_out1_9;

  
  Switch2_out1_2 <= Switch3_out1_6 WHEN Bit_Slice13_out1_2 = '0' ELSE
      Switch3_out1_10;

  Delay_rsvd_4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1_4 <= '0';
      ELSIF enb = '1' THEN
        Delay_out1_4 <= Switch2_out1_2;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_4_process;


  Delay12_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay12_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay12_out1 <= Delay_out1_4;
      END IF;
    END IF;
  END PROCESS Delay12_process;


  BitSlice1_out1 <= mant_a_ext_mant_b_shifted_out1(0);

  sticky_bitget_Sum_1_out1 <= BitSlice1_out1 OR Delay_out1_4;

  Delay4_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1_2 <= '0';
      ELSIF enb = '1' THEN
        Delay4_out1_2 <= sticky_bitget_Sum_1_out1;
      END IF;
    END IF;
  END PROCESS Delay4_2_process;


  
  if_bitget_Sum_Sum_WordLength_2_out1 <= Delay12_out1 WHEN Delay3_out1_1 = '0' ELSE
      Delay4_out1_2;

  BitSlice_out1_1 <= BitSlice6_out1(0);

  BitSlice1_out1_1 <= BitSlice6_out1(1);

  Delay19_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay19_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay19_out1 <= if_bitget_Sum_Sum_WordLength_2_out1;
      END IF;
    END IF;
  END PROCESS Delay19_process;


  sticky_bitget_Sum_1_out1_1 <= BitSlice5_out1 OR Delay19_out1;

  alphabitget_Mant_tmp_2_0_out1 <= BitSlice1_out1_1 OR sticky_bitget_Sum_1_out1_1;

  alphabitget_Mant_tmp_1_0_out1 <= BitSlice_out1_1 AND alphabitget_Mant_tmp_2_0_out1;

  alpha0_out1_2 <= '0';

  BitSlice4_out1 <= BitSlice6_out1(23 DOWNTO 1);

  Bit_Concat_out1_3 <= alpha0_out1_2 & BitSlice4_out1;

  cast_2_like_Mant_tmp_out1 <= to_unsigned(16#000001#, 24);

  Mant_tmp_cast_2_like_Man_out1 <= Bit_Concat_out1_3 + cast_2_like_Mant_tmp_out1;

  
  if_bitget_Mant_tmp_1_0_out1 <= Bit_Concat_out1_3 WHEN alphabitget_Mant_tmp_1_0_out1 = '0' ELSE
      Mant_tmp_cast_2_like_Man_out1;

  BitSlice2_out1 <= if_bitget_Mant_tmp_1_0_out1(23);

  BitSlice4_out1_1 <= Delay15_out1(25);

  C4_out1 <= to_unsigned(16#00#, 8);

  
  Sum_0_out1 <= '1' WHEN Delay1_out1_3 = to_unsigned(16#0000000#, 27) ELSE
      '0';

  exp_a_cor_shift_length_out1 <= Delay2_out1_1 - resize(Delay_out1_3, 8);

  C2_out1 <= to_unsigned(16#01#, 8);

  
  if_shift_length_exp_a_cor_out1 <= exp_a_cor_shift_length_out1 WHEN Logical_Operator1_out1_3 = '0' ELSE
      C2_out1;

  BitSlice2_out1_1 <= Delay1_out1_3(25);

  C3_out1 <= to_unsigned(16#00#, 8);

  
  if_Sum_0_out1 <= if_shift_length_exp_a_cor_out1 WHEN Sum_0_out1 = '0' ELSE
      C3_out1;

  
  if_bitget_Sum_Sum_WordLength_1_out1 <= if_Sum_0_out1 WHEN BitSlice2_out1_1 = '0' ELSE
      Delay2_out1_1;

  C_out1_2 <= to_unsigned(16#01#, 8);

  exp_a_cor_1_out1_1 <= C_out1_2 + Delay2_out1_1;

  
  if_bitget_Sum_Sum_WordLength_1_out1_1 <= if_bitget_Sum_Sum_WordLength_1_out1 WHEN Delay3_out1_1 = '0' ELSE
      exp_a_cor_1_out1_1;

  Delay14_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay14_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay14_out1 <= if_bitget_Sum_Sum_WordLength_1_out1_1;
      END IF;
    END IF;
  END PROCESS Delay14_process;


  
  if_bitget_Sum_Sum_WordLength_out1_1 <= C4_out1 WHEN BitSlice4_out1_1 = '0' ELSE
      Delay14_out1;

  cast_1_like_Exp_out1 <= to_unsigned(16#01#, 8);

  Exp_cast_1_like_Exp_out1 <= if_bitget_Sum_Sum_WordLength_out1_1 + cast_1_like_Exp_out1;

  
  if_bitget_Mant_tmp_Mant_tmp_Wor_out1 <= if_bitget_Sum_Sum_WordLength_out1_1 WHEN BitSlice2_out1 = '0' ELSE
      Exp_cast_1_like_Exp_out1;

  
  Exponent_0_out1_2 <= '1' WHEN if_bitget_Mant_tmp_Mant_tmp_Wor_out1 = to_unsigned(16#00#, 8) ELSE
      '0';

  BitSlice3_out1_1 <= if_bitget_Mant_tmp_1_0_out1(22 DOWNTO 0);

  
  Mantissa_0_out1 <= '1' WHEN BitSlice3_out1_1 = to_unsigned(16#000000#, 23) ELSE
      '0';

  alphaExponent_0_Mantissa_out1 <= Exponent_0_out1_2 AND Mantissa_0_out1;

  Constant_out1_2 <= '0';

  
  Switch_out1_1 <= alphaExponent_0_Mantissa_out1 WHEN Delay18_out1 = '0' ELSE
      Constant_out1_2;

  Delay12_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay12_out1_1 <= '0';
      ELSIF enb = '1' THEN
        Delay12_out1_1 <= if_bitconcat_aExponent_aMantiss_2_ou_1;
      END IF;
    END IF;
  END PROCESS Delay12_1_process;


  Delay29_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay29_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay29_out1 <= Delay12_out1_1;
      END IF;
    END IF;
  END PROCESS Delay29_process;


  Delay14_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay14_reg_rsvd(0) <= '0';
        Delay14_reg_rsvd(1) <= '0';
      ELSIF enb = '1' THEN
        Delay14_reg_rsvd(0) <= Delay14_reg_next(0);
        Delay14_reg_rsvd(1) <= Delay14_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay14_1_process;

  Delay14_out1_1 <= Delay14_reg_rsvd(1);
  Delay14_reg_next(0) <= Delay29_out1;
  Delay14_reg_next(1) <= Delay14_reg_rsvd(0);

  alphaaSign_1_bSign_1_out1 <= if_bitconcat_aExponent_aMantiss_2_ou_1 AND 
    if_bitconcat_aExponent_aMantiss_5_ou_1;

  Delay9_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay9_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay9_out1 <= alphaaSign_1_bSign_1_out1;
      END IF;
    END IF;
  END PROCESS Delay9_process;


  Delay25_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay25_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay25_out1 <= Delay9_out1;
      END IF;
    END IF;
  END PROCESS Delay25_process;


  Delay13_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay13_reg_rsvd(0) <= '0';
        Delay13_reg_rsvd(1) <= '0';
      ELSIF enb = '1' THEN
        Delay13_reg_rsvd(0) <= Delay13_reg_next(0);
        Delay13_reg_rsvd(1) <= Delay13_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay13_1_process;

  Delay13_out1_1 <= Delay13_reg_rsvd(1);
  Delay13_reg_next(0) <= Delay25_out1;
  Delay13_reg_next(1) <= Delay13_reg_rsvd(0);

  
  if_Exponent_0_Mantissa_out1 <= Delay14_out1_1 WHEN Switch_out1_1 = '0' ELSE
      Delay13_out1_1;

  Delay6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay6_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay6_out1 <= if_Exponent_0_Mantissa_out1;
      END IF;
    END IF;
  END PROCESS Delay6_process;


  Delay32_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay32_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay32_out1 <= if_bitconcat_aExponent_aMantiss_out1;
      END IF;
    END IF;
  END PROCESS Delay32_process;


  Delay34_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay34_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay34_out1 <= Delay32_out1;
      END IF;
    END IF;
  END PROCESS Delay34_process;


  Delay15_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay15_reg_rsvd(0) <= to_unsigned(16#00#, 8);
        Delay15_reg_rsvd(1) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay15_reg_rsvd(0) <= Delay15_reg_next(0);
        Delay15_reg_rsvd(1) <= Delay15_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay15_1_process;

  Delay15_out1_1 <= Delay15_reg_rsvd(1);
  Delay15_reg_next(0) <= Delay34_out1;
  Delay15_reg_next(1) <= Delay15_reg_rsvd(0);

  
  if_aExponent_cfType_Exponent_out1 <= if_bitget_Mant_tmp_Mant_tmp_Wor_out1 WHEN Delay18_out1 = '0' ELSE
      Delay15_out1_1;

  Delay7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay7_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay7_out1 <= if_aExponent_cfType_Exponent_out1;
      END IF;
    END IF;
  END PROCESS Delay7_process;


  opp_signs_exp_b_cfType_out1 <= bitxor_out1 AND exp_b_cfType_Exponent_Inf_o_out1;

  
  mant_a_0_out1 <= '1' WHEN if_bitconcat_aExponent_aMantiss_1_ou_1 /= to_unsigned(16#000000#, 23) ELSE
      '0';

  alphamant_a_0_opp_signs_out1 <= opp_signs_exp_b_cfType_out1 OR mant_a_0_out1;

  BitSet_out1 <= if_bitconcat_aExponent_aMantiss_1_ou_1 OR to_unsigned(16#400000#, 23);

  
  if_mant_a_0_opp_signs_out1 <= if_bitconcat_aExponent_aMantiss_1_ou_1 WHEN alphamant_a_0_opp_signs_out1 = 
    '0' ELSE
      BitSet_out1;

  Delay2_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_3 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay2_out1_3 <= if_mant_a_0_opp_signs_out1;
      END IF;
    END IF;
  END PROCESS Delay2_3_process;


  Delay38_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay38_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay38_out1 <= Delay2_out1_3;
      END IF;
    END IF;
  END PROCESS Delay38_process;


  Delay17_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay17_reg_rsvd(0) <= to_unsigned(16#000000#, 23);
        Delay17_reg_rsvd(1) <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay17_reg_rsvd(0) <= Delay17_reg_next(0);
        Delay17_reg_rsvd(1) <= Delay17_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay17_process;

  Delay17_out1 <= Delay17_reg_rsvd(1);
  Delay17_reg_next(0) <= Delay38_out1;
  Delay17_reg_next(1) <= Delay17_reg_rsvd(0);

  
  if_aExponent_cfType_Exponent_1_out1 <= BitSlice3_out1_1 WHEN Delay18_out1 = '0' ELSE
      Delay17_out1;

  Delay8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay8_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay8_out1 <= if_aExponent_cfType_Exponent_1_out1;
      END IF;
    END IF;
  END PROCESS Delay8_process;


  -- Combine FP sign, exponent, mantissa into 32 bit word
  nfp_out_pack <= Delay6_out1 & Delay7_out1 & Delay8_out1;

  nfp_out <= std_logic_vector(nfp_out_pack);

END rtl;

