LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY nfp_mul_single IS
  PORT( clk                               :   IN    std_logic;
        reset_x                           :   IN    std_logic;
        enb                               :   IN    std_logic;
        nfp_in1                           :   IN    std_logic_vector(31 DOWNTO 0);
        nfp_in2                           :   IN    std_logic_vector(31 DOWNTO 0);
        nfp_out                           :   OUT   std_logic_vector(31 DOWNTO 0)
        );
END nfp_mul_single;


ARCHITECTURE rtl OF nfp_mul_single IS

  -- Signals
  SIGNAL nfp_in2_unsigned                 : unsigned(31 DOWNTO 0);
  SIGNAL BS                               : std_logic;
  SIGNAL BE                               : unsigned(7 DOWNTO 0);
  SIGNAL BM                               : unsigned(22 DOWNTO 0);
  SIGNAL Compare_To_Constant1_out1        : std_logic;
  SIGNAL Delay16_out1                     : std_logic;
  SIGNAL Compare_To_Zero3_out1            : std_logic;
  SIGNAL Delay14_out1                     : std_logic;
  SIGNAL Logical_Operator1_out1           : std_logic;
  SIGNAL nfp_in1_unsigned                 : unsigned(31 DOWNTO 0);
  SIGNAL AS                               : std_logic;
  SIGNAL AE                               : unsigned(7 DOWNTO 0);
  SIGNAL AM                               : unsigned(22 DOWNTO 0);
  SIGNAL Compare_To_Constant_out1         : std_logic;
  SIGNAL Delay21_out1                     : std_logic;
  SIGNAL Compare_To_Zero2_out1            : std_logic;
  SIGNAL Delay19_out1                     : std_logic;
  SIGNAL Logical_Operator_out1            : std_logic;
  SIGNAL Delay3_out1                      : std_logic;
  SIGNAL Delay7_out1                      : std_logic;
  SIGNAL Logical_Operator_out1_1          : std_logic;
  SIGNAL Switch_out1                      : std_logic;
  SIGNAL Switch1_out1                     : std_logic;
  SIGNAL Delay29_reg_rsvd                 : std_logic_vector(0 TO 2);
  SIGNAL Delay29_reg_next                 : std_logic_vector(0 TO 2);
  SIGNAL Delay29_out1                     : std_logic;
  SIGNAL Delay_reg_rsvd                   : std_logic_vector(0 TO 1);
  SIGNAL Delay_reg_next                   : std_logic_vector(0 TO 1);
  SIGNAL Delay_out1                       : std_logic;
  SIGNAL Constant8_out1                   : std_logic;
  SIGNAL Constant7_out1                   : unsigned(7 DOWNTO 0);
  SIGNAL Relational_Operator_relop1       : std_logic;
  SIGNAL Delay4_out1                      : std_logic;
  SIGNAL Logical_Operator2_out1           : std_logic;
  SIGNAL Logical_Operator_out1_2          : std_logic;
  SIGNAL Add_out1                         : unsigned(7 DOWNTO 0);
  SIGNAL Delay3_out1_1                    : unsigned(7 DOWNTO 0);
  SIGNAL Add_add_cast                     : unsigned(7 DOWNTO 0);
  SIGNAL Constant6_out1                   : unsigned(7 DOWNTO 0);
  SIGNAL Compare_To_Zero_out1             : std_logic;
  SIGNAL Delay23_out1                     : std_logic;
  SIGNAL Constant1_out1                   : std_logic;
  SIGNAL Constant_out1                    : std_logic;
  SIGNAL Switch1_out1_1                   : std_logic;
  SIGNAL Delay6_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Concat_out1                  : unsigned(23 DOWNTO 0);
  SIGNAL Constant5_out1                   : unsigned(23 DOWNTO 0);
  SIGNAL Switch_out1_1                    : unsigned(23 DOWNTO 0);
  SIGNAL Delay2_out1                      : unsigned(23 DOWNTO 0);
  SIGNAL Logical_Operator3_out1           : std_logic;
  SIGNAL Compare_To_Zero1_out1            : std_logic;
  SIGNAL Delay20_out1                     : std_logic;
  SIGNAL Constant3_out1                   : std_logic;
  SIGNAL Constant2_out1                   : std_logic;
  SIGNAL Switch2_out1                     : std_logic;
  SIGNAL Logical_Operator_out1_3          : std_logic;
  SIGNAL Delay8_out1                      : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Concat1_out1                 : unsigned(23 DOWNTO 0);
  SIGNAL Constant4_out1                   : unsigned(23 DOWNTO 0);
  SIGNAL Switch3_out1                     : unsigned(23 DOWNTO 0);
  SIGNAL Delay1_out1                      : unsigned(23 DOWNTO 0);
  SIGNAL Product_out1                     : unsigned(47 DOWNTO 0);
  SIGNAL Delay4_out1_1                    : unsigned(47 DOWNTO 0);
  SIGNAL Constant1_out1_1                 : std_logic;
  SIGNAL Bit_Concat_out1_1                : unsigned(48 DOWNTO 0);
  SIGNAL Compare_To_Zero1_out1_1          : std_logic;
  SIGNAL Logical_Operator1_out1_1         : std_logic;
  SIGNAL Delay4_out1_2                    : unsigned(7 DOWNTO 0);
  SIGNAL Delay5_out1                      : unsigned(7 DOWNTO 0);
  SIGNAL Subtract_out1                    : unsigned(8 DOWNTO 0);
  SIGNAL Delay_out1_1                     : unsigned(8 DOWNTO 0);
  SIGNAL Constant2_out1_1                 : unsigned(6 DOWNTO 0);
  SIGNAL Constant1_out1_2                 : std_logic;
  SIGNAL Constant3_out1_1                 : std_logic;
  SIGNAL Switch_out1_2                    : std_logic;
  SIGNAL Bit_Concat1_out1_1               : unsigned(7 DOWNTO 0);
  SIGNAL Switch1_out1_2                   : std_logic;
  SIGNAL Bit_Concat_out1_2                : unsigned(7 DOWNTO 0);
  SIGNAL Add1_out1                        : unsigned(8 DOWNTO 0);
  SIGNAL Delay3_out1_2                    : std_logic;
  SIGNAL Delay2_out1_1                    : unsigned(8 DOWNTO 0);
  SIGNAL Subtract2_sub_cast               : signed(31 DOWNTO 0);
  SIGNAL Subtract2_sub_cast_1             : signed(31 DOWNTO 0);
  SIGNAL Subtract2_sub_temp               : signed(31 DOWNTO 0);
  SIGNAL Subtract2_out1                   : signed(9 DOWNTO 0);
  SIGNAL Constant4_out1_1                 : signed(9 DOWNTO 0);
  SIGNAL Switch2_out1_1                   : signed(9 DOWNTO 0);
  SIGNAL Delay27_out1                     : signed(9 DOWNTO 0);
  SIGNAL Constant_out1_1                  : signed(9 DOWNTO 0);
  SIGNAL Switch1_out1_3                   : signed(9 DOWNTO 0);
  SIGNAL Delay5_out1_1                    : signed(9 DOWNTO 0);
  SIGNAL Bit_Slice25_out1                 : std_logic;
  SIGNAL Constant25_out1                  : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice24_out1                 : std_logic;
  SIGNAL Constant24_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch24_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice23_out1                 : std_logic;
  SIGNAL Constant23_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch23_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice22_out1                 : std_logic;
  SIGNAL Constant22_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch22_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice21_out1                 : std_logic;
  SIGNAL Constant21_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch21_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice10_out1                 : std_logic;
  SIGNAL Constant20_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch20_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice19_out1                 : std_logic;
  SIGNAL Constant19_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch19_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice18_out1                 : std_logic;
  SIGNAL Constant18_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch18_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice17_out1                 : std_logic;
  SIGNAL Constant17_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch17_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice16_out1                 : std_logic;
  SIGNAL Constant16_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch16_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice15_out1                 : std_logic;
  SIGNAL Constant15_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch15_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice14_out1                 : std_logic;
  SIGNAL Constant14_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch14_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice13_out1                 : std_logic;
  SIGNAL Constant13_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch13_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice12_out1                 : std_logic;
  SIGNAL Constant12_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch12_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice11_out1                 : std_logic;
  SIGNAL Constant11_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch11_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice_out1                   : std_logic;
  SIGNAL Constant10_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch10_out1                    : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice9_out1                  : std_logic;
  SIGNAL Constant9_out1                   : signed(5 DOWNTO 0);
  SIGNAL Switch9_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice8_out1                  : std_logic;
  SIGNAL Constant8_out1_1                 : signed(5 DOWNTO 0);
  SIGNAL Switch8_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice7_out1                  : std_logic;
  SIGNAL Constant7_out1_1                 : signed(5 DOWNTO 0);
  SIGNAL Switch7_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice6_out1                  : std_logic;
  SIGNAL Constant6_out1_1                 : signed(5 DOWNTO 0);
  SIGNAL Switch6_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice5_out1                  : std_logic;
  SIGNAL Constant5_out1_1                 : signed(5 DOWNTO 0);
  SIGNAL Switch5_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice4_out1                  : std_logic;
  SIGNAL Constant4_out1_2                 : signed(5 DOWNTO 0);
  SIGNAL Switch4_out1                     : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice3_out1                  : std_logic;
  SIGNAL Constant3_out1_2                 : signed(5 DOWNTO 0);
  SIGNAL Switch3_out1_1                   : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice2_out1                  : std_logic;
  SIGNAL Constant2_out1_2                 : signed(5 DOWNTO 0);
  SIGNAL Switch2_out1_2                   : signed(5 DOWNTO 0);
  SIGNAL Bit_Slice1_out1                  : std_logic;
  SIGNAL Constant1_out1_3                 : signed(5 DOWNTO 0);
  SIGNAL Switch1_out1_4                   : signed(5 DOWNTO 0);
  SIGNAL Constant26_out1                  : signed(5 DOWNTO 0);
  SIGNAL Switch_out1_3                    : signed(5 DOWNTO 0);
  SIGNAL Delay1_out1_1                    : signed(5 DOWNTO 0);
  SIGNAL Add_sub_temp                     : signed(31 DOWNTO 0);
  SIGNAL Add_out1_1                       : signed(9 DOWNTO 0);
  SIGNAL Compare_To_Constant_out1_1       : std_logic;
  SIGNAL Constant1_out1_4                 : signed(8 DOWNTO 0);
  SIGNAL Constant1_out1_dtc               : signed(9 DOWNTO 0);
  SIGNAL Switch_out1_4                    : signed(9 DOWNTO 0);
  SIGNAL Delay18_out1                     : signed(9 DOWNTO 0);
  SIGNAL Compare_To_Constant1_out1_1      : std_logic;
  SIGNAL Logical_Operator1_out1_2         : std_logic;
  SIGNAL Logical_Operator4_out1           : std_logic;
  SIGNAL Logical_Operator7_out1           : std_logic;
  SIGNAL Logical_Operator5_out1           : std_logic;
  SIGNAL Logical_Operator6_out1           : std_logic;
  SIGNAL Logical_Operator8_out1           : std_logic;
  SIGNAL Inf_Zero_out1                    : std_logic;
  SIGNAL Logical_Operator2_out1_1         : std_logic;
  SIGNAL Logical_Operator10_out1          : std_logic;
  SIGNAL Delay22_reg_rsvd                 : std_logic_vector(0 TO 2);
  SIGNAL Delay22_reg_next                 : std_logic_vector(0 TO 2);
  SIGNAL Delay22_out1                     : std_logic;
  SIGNAL Delay13_out1                     : std_logic;
  SIGNAL Logical_Operator_out1_4          : std_logic;
  SIGNAL Compare_To_Constant_out1_2       : std_logic;
  SIGNAL Constant1_out1_5                 : unsigned(7 DOWNTO 0);
  SIGNAL Delay2_out1_2                    : unsigned(48 DOWNTO 0);
  SIGNAL Compare_To_Zero_out1_1           : std_logic;
  SIGNAL Bit_Slice_out1_1                 : unsigned(4 DOWNTO 0);
  SIGNAL Shift_Arithmetic_out1            : unsigned(48 DOWNTO 0);
  SIGNAL Bit_Shift_out1                   : unsigned(48 DOWNTO 0);
  SIGNAL Delay3_out1_3                    : unsigned(48 DOWNTO 0);
  SIGNAL Switch_out1_5                    : unsigned(48 DOWNTO 0);
  SIGNAL Constant_out1_2                  : signed(8 DOWNTO 0);
  SIGNAL Subtract_sub_temp                : signed(31 DOWNTO 0);
  SIGNAL Subtract_out1_1                  : signed(15 DOWNTO 0);
  SIGNAL Compare_To_Constant_out1_3       : std_logic;
  SIGNAL Subtract_out1_dtc                : signed(5 DOWNTO 0);
  SIGNAL Compare_To_Constant1_out1_2      : std_logic;
  SIGNAL Constant1_out1_6                 : signed(5 DOWNTO 0);
  SIGNAL Switch_out1_6                    : signed(5 DOWNTO 0);
  SIGNAL Constant2_out1_3                 : signed(5 DOWNTO 0);
  SIGNAL Switch1_out1_5                   : signed(5 DOWNTO 0);
  SIGNAL Unary_Minus_in0                  : signed(6 DOWNTO 0);
  SIGNAL Unary_Minus_out1                 : signed(5 DOWNTO 0);
  SIGNAL shift_arithmetic_shift_direction : std_logic;
  SIGNAL Constant_out1_3                  : unsigned(30 DOWNTO 0);
  SIGNAL Bit_Concat_out1_3                : unsigned(79 DOWNTO 0);
  SIGNAL shift_arithmetic_abs_y           : signed(6 DOWNTO 0);
  SIGNAL shift_arithmetic_shift_value     : unsigned(6 DOWNTO 0);
  SIGNAL shift_arithmetic_right           : unsigned(79 DOWNTO 0);
  SIGNAL shift_arithmetic_left            : unsigned(79 DOWNTO 0);
  SIGNAL Shift_Arithmetic_out1_1          : unsigned(79 DOWNTO 0);
  SIGNAL Bit_Slice1_out1_1                : unsigned(30 DOWNTO 0);
  SIGNAL Bit_Slice_out1_2                 : unsigned(48 DOWNTO 0);
  SIGNAL Bit_Set_out1                     : unsigned(48 DOWNTO 0);
  SIGNAL Switch2_out1_3                   : unsigned(48 DOWNTO 0);
  SIGNAL Switch1_out1_6                   : unsigned(48 DOWNTO 0);
  SIGNAL Bit_Slice_out1_3                 : unsigned(47 DOWNTO 0);
  SIGNAL Bit_Slice2_out1_1                : unsigned(1 DOWNTO 0);
  SIGNAL Bit_Slice4_out1_1                : std_logic;
  SIGNAL Bit_Slice1_out1_2                : unsigned(21 DOWNTO 0);
  SIGNAL Bit_Reduce_out1                  : std_logic;
  SIGNAL Bit_Slice5_out1_1                : std_logic;
  SIGNAL Bit_Slice3_out1_1                : std_logic;
  SIGNAL Logical_Operator1_out1_3         : std_logic;
  SIGNAL Logical_Operator_out1_5          : std_logic;
  SIGNAL Delay1_out1_2                    : std_logic;
  SIGNAL Bit_Slice1_out1_3                : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Slice1_out1_4                : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Slice1_out1_dtc              : unsigned(23 DOWNTO 0);
  SIGNAL Constant_out1_4                  : std_logic;
  SIGNAL Add_add_cast_1                   : unsigned(31 DOWNTO 0);
  SIGNAL Add_out1_2                       : unsigned(23 DOWNTO 0);
  SIGNAL Switch_out1_7                    : unsigned(23 DOWNTO 0);
  SIGNAL Bit_Slice2_out1_2                : std_logic;
  SIGNAL Add1_add_cast                    : unsigned(31 DOWNTO 0);
  SIGNAL Add1_out1_1                      : unsigned(7 DOWNTO 0);
  SIGNAL Add_add_cast_2                   : signed(31 DOWNTO 0);
  SIGNAL Add_add_temp                     : signed(31 DOWNTO 0);
  SIGNAL Add_out1_3                       : unsigned(7 DOWNTO 0);
  SIGNAL Constant1_out1_7                 : unsigned(7 DOWNTO 0);
  SIGNAL Switch1_out1_7                   : unsigned(7 DOWNTO 0);
  SIGNAL Constant4_out1_3                 : unsigned(7 DOWNTO 0);
  SIGNAL Switch4_out1_1                   : unsigned(7 DOWNTO 0);
  SIGNAL Switch6_out1_1                   : unsigned(7 DOWNTO 0);
  SIGNAL Delay1_out1_3                    : unsigned(7 DOWNTO 0);
  SIGNAL Bit_Slice4_out1_2                : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Shift_out1_1                 : unsigned(22 DOWNTO 0);
  SIGNAL Switch1_out1_8                   : unsigned(22 DOWNTO 0);
  SIGNAL Constant2_out1_4                 : unsigned(22 DOWNTO 0);
  SIGNAL Switch2_out1_4                   : unsigned(22 DOWNTO 0);
  SIGNAL Constant5_out1_2                 : unsigned(22 DOWNTO 0);
  SIGNAL Bit_Set_out1_1                   : unsigned(22 DOWNTO 0);
  SIGNAL Switch7_out1_1                   : unsigned(22 DOWNTO 0);
  SIGNAL Switch5_out1_1                   : unsigned(22 DOWNTO 0);
  SIGNAL Delay2_out1_3                    : unsigned(22 DOWNTO 0);
  SIGNAL nfp_out_pack                     : unsigned(31 DOWNTO 0);

BEGIN
  nfp_in2_unsigned <= unsigned(nfp_in2);

  -- Split 32 bit word into FP sign, exponent, mantissa
  BS <= nfp_in2_unsigned(31);
  BE <= nfp_in2_unsigned(30 DOWNTO 23);
  BM <= nfp_in2_unsigned(22 DOWNTO 0);

  
  Compare_To_Constant1_out1 <= '1' WHEN BE = to_unsigned(16#FF#, 8) ELSE
      '0';

  Delay16_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay16_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay16_out1 <= Compare_To_Constant1_out1;
      END IF;
    END IF;
  END PROCESS Delay16_process;


  
  Compare_To_Zero3_out1 <= '1' WHEN BM /= to_unsigned(16#000000#, 23) ELSE
      '0';

  Delay14_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay14_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay14_out1 <= Compare_To_Zero3_out1;
      END IF;
    END IF;
  END PROCESS Delay14_process;


  Logical_Operator1_out1 <= Delay16_out1 AND Delay14_out1;

  nfp_in1_unsigned <= unsigned(nfp_in1);

  -- Split 32 bit word into FP sign, exponent, mantissa
  AS <= nfp_in1_unsigned(31);
  AE <= nfp_in1_unsigned(30 DOWNTO 23);
  AM <= nfp_in1_unsigned(22 DOWNTO 0);

  
  Compare_To_Constant_out1 <= '1' WHEN AE = to_unsigned(16#FF#, 8) ELSE
      '0';

  Delay21_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay21_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay21_out1 <= Compare_To_Constant_out1;
      END IF;
    END IF;
  END PROCESS Delay21_process;


  
  Compare_To_Zero2_out1 <= '1' WHEN AM /= to_unsigned(16#000000#, 23) ELSE
      '0';

  Delay19_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay19_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay19_out1 <= Compare_To_Zero2_out1;
      END IF;
    END IF;
  END PROCESS Delay19_process;


  Logical_Operator_out1 <= Delay21_out1 AND Delay19_out1;

  Delay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay3_out1 <= AS;
      END IF;
    END IF;
  END PROCESS Delay3_process;


  Delay7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay7_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay7_out1 <= BS;
      END IF;
    END IF;
  END PROCESS Delay7_process;


  Logical_Operator_out1_1 <= Delay3_out1 XOR Delay7_out1;

  
  Switch_out1 <= Logical_Operator_out1_1 WHEN Logical_Operator_out1 = '0' ELSE
      Delay3_out1;

  
  Switch1_out1 <= Switch_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Delay7_out1;

  Delay29_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay29_reg_rsvd(0) <= '0';
        Delay29_reg_rsvd(1) <= '0';
        Delay29_reg_rsvd(2) <= '0';
      ELSIF enb = '1' THEN
        Delay29_reg_rsvd(0) <= Delay29_reg_next(0);
        Delay29_reg_rsvd(1) <= Delay29_reg_next(1);
        Delay29_reg_rsvd(2) <= Delay29_reg_next(2);
      END IF;
    END IF;
  END PROCESS Delay29_process;

  Delay29_out1 <= Delay29_reg_rsvd(2);
  Delay29_reg_next(0) <= Switch1_out1;
  Delay29_reg_next(1) <= Delay29_reg_rsvd(0);
  Delay29_reg_next(2) <= Delay29_reg_rsvd(1);

  Delay_rsvd_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_reg_rsvd(0) <= '0';
        Delay_reg_rsvd(1) <= '0';
      ELSIF enb = '1' THEN
        Delay_reg_rsvd(0) <= Delay_reg_next(0);
        Delay_reg_rsvd(1) <= Delay_reg_next(1);
      END IF;
    END IF;
  END PROCESS Delay_rsvd_process;

  Delay_out1 <= Delay_reg_rsvd(1);
  Delay_reg_next(0) <= Delay29_out1;
  Delay_reg_next(1) <= Delay_reg_rsvd(0);

  Constant8_out1 <= '1';

  Constant7_out1 <= to_unsigned(16#06#, 8);

  Delay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay4_out1 <= Relational_Operator_relop1;
      END IF;
    END IF;
  END PROCESS Delay4_process;


  Logical_Operator2_out1 <=  NOT Delay4_out1;

  Logical_Operator_out1_2 <= Constant8_out1 AND Logical_Operator2_out1;

  Delay3_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay3_out1_1 <= Add_out1;
      END IF;
    END IF;
  END PROCESS Delay3_1_process;


  Add_add_cast <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & Logical_Operator_out1_2;
  Add_out1 <= Delay3_out1_1 + Add_add_cast;

  
  Relational_Operator_relop1 <= '1' WHEN Add_out1 >= Constant7_out1 ELSE
      '0';

  Constant6_out1 <= to_unsigned(16#00#, 8);

  
  Compare_To_Zero_out1 <= '1' WHEN AE = to_unsigned(16#00#, 8) ELSE
      '0';

  Delay23_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay23_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay23_out1 <= Compare_To_Zero_out1;
      END IF;
    END IF;
  END PROCESS Delay23_process;


  Constant1_out1 <= '1';

  Constant_out1 <= '0';

  
  Switch1_out1_1 <= Constant1_out1 WHEN Delay23_out1 = '0' ELSE
      Constant_out1;

  Delay6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay6_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay6_out1 <= AM;
      END IF;
    END IF;
  END PROCESS Delay6_process;


  Bit_Concat_out1 <= Switch1_out1_1 & Delay6_out1;

  Constant5_out1 <= to_unsigned(16#800000#, 24);

  
  Switch_out1_1 <= Bit_Concat_out1 WHEN Logical_Operator1_out1 = '0' ELSE
      Constant5_out1;

  Delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1 <= to_unsigned(16#000000#, 24);
      ELSIF enb = '1' THEN
        Delay2_out1 <= Switch_out1_1;
      END IF;
    END IF;
  END PROCESS Delay2_process;


  Logical_Operator3_out1 <=  NOT Logical_Operator1_out1;

  
  Compare_To_Zero1_out1 <= '1' WHEN BE = to_unsigned(16#00#, 8) ELSE
      '0';

  Delay20_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay20_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay20_out1 <= Compare_To_Zero1_out1;
      END IF;
    END IF;
  END PROCESS Delay20_process;


  Constant3_out1 <= '1';

  Constant2_out1 <= '0';

  
  Switch2_out1 <= Constant3_out1 WHEN Delay20_out1 = '0' ELSE
      Constant2_out1;

  Logical_Operator_out1_3 <= Logical_Operator_out1 AND Logical_Operator3_out1;

  Delay8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay8_out1 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay8_out1 <= BM;
      END IF;
    END IF;
  END PROCESS Delay8_process;


  Bit_Concat1_out1 <= Switch2_out1 & Delay8_out1;

  Constant4_out1 <= to_unsigned(16#800000#, 24);

  
  Switch3_out1 <= Bit_Concat1_out1 WHEN Logical_Operator_out1_3 = '0' ELSE
      Constant4_out1;

  Delay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1 <= to_unsigned(16#000000#, 24);
      ELSIF enb = '1' THEN
        Delay1_out1 <= Switch3_out1;
      END IF;
    END IF;
  END PROCESS Delay1_process;


  Product_out1 <= Delay2_out1 * Delay1_out1;

  Delay4_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1_1 <= to_unsigned(0, 48);
      ELSIF enb = '1' THEN
        Delay4_out1_1 <= Product_out1;
      END IF;
    END IF;
  END PROCESS Delay4_1_process;


  Constant1_out1_1 <= '0';

  Bit_Concat_out1_1 <= Delay4_out1_1 & Constant1_out1_1;

  
  Compare_To_Zero1_out1_1 <= '1' WHEN Bit_Concat_out1_1 = to_unsigned(0, 49) ELSE
      '0';

  Logical_Operator1_out1_1 <= Delay21_out1 OR Delay16_out1;

  Delay4_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay4_out1_2 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay4_out1_2 <= AE;
      END IF;
    END IF;
  END PROCESS Delay4_2_process;


  Delay5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay5_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay5_out1 <= BE;
      END IF;
    END IF;
  END PROCESS Delay5_process;


  Subtract_out1 <= resize(resize(Delay4_out1_2, 32) + resize(Delay5_out1, 32), 9);

  Delay_rsvd_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay_out1_1 <= to_unsigned(16#000#, 9);
      ELSIF enb = '1' THEN
        Delay_out1_1 <= Subtract_out1;
      END IF;
    END IF;
  END PROCESS Delay_rsvd_1_process;


  Constant2_out1_1 <= to_unsigned(16#3F#, 7);

  Constant1_out1_2 <= '1';

  Constant3_out1_1 <= '0';

  
  Switch_out1_2 <= Constant1_out1_2 WHEN Delay23_out1 = '0' ELSE
      Constant3_out1_1;

  Bit_Concat1_out1_1 <= Constant2_out1_1 & Switch_out1_2;

  
  Switch1_out1_2 <= Constant1_out1_2 WHEN Delay20_out1 = '0' ELSE
      Constant3_out1_1;

  Bit_Concat_out1_2 <= Constant2_out1_1 & Switch1_out1_2;

  Add1_out1 <= resize(resize(Bit_Concat1_out1_1, 32) + resize(Bit_Concat_out1_2, 32), 9);

  Delay3_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1_2 <= '0';
      ELSIF enb = '1' THEN
        Delay3_out1_2 <= Logical_Operator1_out1_1;
      END IF;
    END IF;
  END PROCESS Delay3_2_process;


  Delay2_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_1 <= to_unsigned(16#000#, 9);
      ELSIF enb = '1' THEN
        Delay2_out1_1 <= Add1_out1;
      END IF;
    END IF;
  END PROCESS Delay2_1_process;


  Subtract2_sub_cast <= signed(resize(Delay_out1_1, 32));
  Subtract2_sub_cast_1 <= signed(resize(Delay2_out1_1, 32));
  Subtract2_sub_temp <= Subtract2_sub_cast - Subtract2_sub_cast_1;
  Subtract2_out1 <= Subtract2_sub_temp(9 DOWNTO 0);

  Constant4_out1_1 <= to_signed(16#0FF#, 10);

  
  Switch2_out1_1 <= Subtract2_out1 WHEN Delay3_out1_2 = '0' ELSE
      Constant4_out1_1;

  Delay27_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay27_out1 <= to_signed(16#000#, 10);
      ELSIF enb = '1' THEN
        Delay27_out1 <= Switch2_out1_1;
      END IF;
    END IF;
  END PROCESS Delay27_process;


  Constant_out1_1 <= to_signed(-16#0FF#, 10);

  
  Switch1_out1_3 <= Delay27_out1 WHEN Compare_To_Zero1_out1_1 = '0' ELSE
      Constant_out1_1;

  Delay5_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay5_out1_1 <= to_signed(16#000#, 10);
      ELSIF enb = '1' THEN
        Delay5_out1_1 <= Switch1_out1_3;
      END IF;
    END IF;
  END PROCESS Delay5_1_process;


  Bit_Slice25_out1 <= Bit_Concat_out1_1(24);

  Constant25_out1 <= to_signed(16#18#, 6);

  Bit_Slice24_out1 <= Bit_Concat_out1_1(25);

  Constant24_out1 <= to_signed(16#17#, 6);

  
  Switch24_out1 <= Constant25_out1 WHEN Bit_Slice25_out1 = '0' ELSE
      Constant24_out1;

  Bit_Slice23_out1 <= Bit_Concat_out1_1(26);

  Constant23_out1 <= to_signed(16#16#, 6);

  
  Switch23_out1 <= Switch24_out1 WHEN Bit_Slice24_out1 = '0' ELSE
      Constant23_out1;

  Bit_Slice22_out1 <= Bit_Concat_out1_1(27);

  Constant22_out1 <= to_signed(16#15#, 6);

  
  Switch22_out1 <= Switch23_out1 WHEN Bit_Slice23_out1 = '0' ELSE
      Constant22_out1;

  Bit_Slice21_out1 <= Bit_Concat_out1_1(28);

  Constant21_out1 <= to_signed(16#14#, 6);

  
  Switch21_out1 <= Switch22_out1 WHEN Bit_Slice22_out1 = '0' ELSE
      Constant21_out1;

  Bit_Slice10_out1 <= Bit_Concat_out1_1(29);

  Constant20_out1 <= to_signed(16#13#, 6);

  
  Switch20_out1 <= Switch21_out1 WHEN Bit_Slice21_out1 = '0' ELSE
      Constant20_out1;

  Bit_Slice19_out1 <= Bit_Concat_out1_1(30);

  Constant19_out1 <= to_signed(16#12#, 6);

  
  Switch19_out1 <= Switch20_out1 WHEN Bit_Slice10_out1 = '0' ELSE
      Constant19_out1;

  Bit_Slice18_out1 <= Bit_Concat_out1_1(31);

  Constant18_out1 <= to_signed(16#11#, 6);

  
  Switch18_out1 <= Switch19_out1 WHEN Bit_Slice19_out1 = '0' ELSE
      Constant18_out1;

  Bit_Slice17_out1 <= Bit_Concat_out1_1(32);

  Constant17_out1 <= to_signed(16#10#, 6);

  
  Switch17_out1 <= Switch18_out1 WHEN Bit_Slice18_out1 = '0' ELSE
      Constant17_out1;

  Bit_Slice16_out1 <= Bit_Concat_out1_1(33);

  Constant16_out1 <= to_signed(16#0F#, 6);

  
  Switch16_out1 <= Switch17_out1 WHEN Bit_Slice17_out1 = '0' ELSE
      Constant16_out1;

  Bit_Slice15_out1 <= Bit_Concat_out1_1(34);

  Constant15_out1 <= to_signed(16#0E#, 6);

  
  Switch15_out1 <= Switch16_out1 WHEN Bit_Slice16_out1 = '0' ELSE
      Constant15_out1;

  Bit_Slice14_out1 <= Bit_Concat_out1_1(35);

  Constant14_out1 <= to_signed(16#0D#, 6);

  
  Switch14_out1 <= Switch15_out1 WHEN Bit_Slice15_out1 = '0' ELSE
      Constant14_out1;

  Bit_Slice13_out1 <= Bit_Concat_out1_1(36);

  Constant13_out1 <= to_signed(16#0C#, 6);

  
  Switch13_out1 <= Switch14_out1 WHEN Bit_Slice14_out1 = '0' ELSE
      Constant13_out1;

  Bit_Slice12_out1 <= Bit_Concat_out1_1(37);

  Constant12_out1 <= to_signed(16#0B#, 6);

  
  Switch12_out1 <= Switch13_out1 WHEN Bit_Slice13_out1 = '0' ELSE
      Constant12_out1;

  Bit_Slice11_out1 <= Bit_Concat_out1_1(38);

  Constant11_out1 <= to_signed(16#0A#, 6);

  
  Switch11_out1 <= Switch12_out1 WHEN Bit_Slice12_out1 = '0' ELSE
      Constant11_out1;

  Bit_Slice_out1 <= Bit_Concat_out1_1(39);

  Constant10_out1 <= to_signed(16#09#, 6);

  
  Switch10_out1 <= Switch11_out1 WHEN Bit_Slice11_out1 = '0' ELSE
      Constant10_out1;

  Bit_Slice9_out1 <= Bit_Concat_out1_1(40);

  Constant9_out1 <= to_signed(16#08#, 6);

  
  Switch9_out1 <= Switch10_out1 WHEN Bit_Slice_out1 = '0' ELSE
      Constant9_out1;

  Bit_Slice8_out1 <= Bit_Concat_out1_1(41);

  Constant8_out1_1 <= to_signed(16#07#, 6);

  
  Switch8_out1 <= Switch9_out1 WHEN Bit_Slice9_out1 = '0' ELSE
      Constant8_out1_1;

  Bit_Slice7_out1 <= Bit_Concat_out1_1(42);

  Constant7_out1_1 <= to_signed(16#06#, 6);

  
  Switch7_out1 <= Switch8_out1 WHEN Bit_Slice8_out1 = '0' ELSE
      Constant7_out1_1;

  Bit_Slice6_out1 <= Bit_Concat_out1_1(43);

  Constant6_out1_1 <= to_signed(16#05#, 6);

  
  Switch6_out1 <= Switch7_out1 WHEN Bit_Slice7_out1 = '0' ELSE
      Constant6_out1_1;

  Bit_Slice5_out1 <= Bit_Concat_out1_1(44);

  Constant5_out1_1 <= to_signed(16#04#, 6);

  
  Switch5_out1 <= Switch6_out1 WHEN Bit_Slice6_out1 = '0' ELSE
      Constant5_out1_1;

  Bit_Slice4_out1 <= Bit_Concat_out1_1(45);

  Constant4_out1_2 <= to_signed(16#03#, 6);

  
  Switch4_out1 <= Switch5_out1 WHEN Bit_Slice5_out1 = '0' ELSE
      Constant4_out1_2;

  Bit_Slice3_out1 <= Bit_Concat_out1_1(46);

  Constant3_out1_2 <= to_signed(16#02#, 6);

  
  Switch3_out1_1 <= Switch4_out1 WHEN Bit_Slice4_out1 = '0' ELSE
      Constant3_out1_2;

  Bit_Slice2_out1 <= Bit_Concat_out1_1(47);

  Constant2_out1_2 <= to_signed(16#01#, 6);

  
  Switch2_out1_2 <= Switch3_out1_1 WHEN Bit_Slice3_out1 = '0' ELSE
      Constant2_out1_2;

  Bit_Slice1_out1 <= Bit_Concat_out1_1(48);

  Constant1_out1_3 <= to_signed(16#00#, 6);

  
  Switch1_out1_4 <= Switch2_out1_2 WHEN Bit_Slice2_out1 = '0' ELSE
      Constant1_out1_3;

  Constant26_out1 <= to_signed(-16#01#, 6);

  
  Switch_out1_3 <= Switch1_out1_4 WHEN Bit_Slice1_out1 = '0' ELSE
      Constant26_out1;

  Delay1_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_1 <= to_signed(16#00#, 6);
      ELSIF enb = '1' THEN
        Delay1_out1_1 <= Switch_out1_3;
      END IF;
    END IF;
  END PROCESS Delay1_1_process;


  Add_sub_temp <= resize(Delay5_out1_1, 32) - resize(Delay1_out1_1, 32);
  Add_out1_1 <= Add_sub_temp(9 DOWNTO 0);

  
  Compare_To_Constant_out1_1 <= '1' WHEN Add_out1_1 <= to_signed(-16#07F#, 10) ELSE
      '0';

  Constant1_out1_4 <= to_signed(-16#07F#, 9);

  Constant1_out1_dtc <= resize(Constant1_out1_4, 10);

  
  Switch_out1_4 <= Add_out1_1 WHEN Compare_To_Constant_out1_1 = '0' ELSE
      Constant1_out1_dtc;

  Delay18_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay18_out1 <= to_signed(16#000#, 10);
      ELSIF enb = '1' THEN
        Delay18_out1 <= Switch_out1_4;
      END IF;
    END IF;
  END PROCESS Delay18_process;


  
  Compare_To_Constant1_out1_1 <= '1' WHEN Delay18_out1 > to_signed(16#07F#, 10) ELSE
      '0';

  Logical_Operator1_out1_2 <=  NOT Delay14_out1;

  Logical_Operator4_out1 <= Logical_Operator1_out1_2 AND Delay20_out1;

  Logical_Operator7_out1 <= Logical_Operator4_out1 AND Delay21_out1;

  Logical_Operator5_out1 <=  NOT Delay19_out1;

  Logical_Operator6_out1 <= Logical_Operator5_out1 AND Delay23_out1;

  Logical_Operator8_out1 <= Logical_Operator6_out1 AND Delay16_out1;

  Inf_Zero_out1 <= Logical_Operator7_out1 OR Logical_Operator8_out1;

  Logical_Operator2_out1_1 <= Logical_Operator_out1 OR Logical_Operator1_out1;

  Logical_Operator10_out1 <= Inf_Zero_out1 OR Logical_Operator2_out1_1;

  Delay22_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay22_reg_rsvd(0) <= '0';
        Delay22_reg_rsvd(1) <= '0';
        Delay22_reg_rsvd(2) <= '0';
      ELSIF enb = '1' THEN
        Delay22_reg_rsvd(0) <= Delay22_reg_next(0);
        Delay22_reg_rsvd(1) <= Delay22_reg_next(1);
        Delay22_reg_rsvd(2) <= Delay22_reg_next(2);
      END IF;
    END IF;
  END PROCESS Delay22_process;

  Delay22_out1 <= Delay22_reg_rsvd(2);
  Delay22_reg_next(0) <= Logical_Operator10_out1;
  Delay22_reg_next(1) <= Delay22_reg_rsvd(0);
  Delay22_reg_next(2) <= Delay22_reg_rsvd(1);

  Delay13_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay13_out1 <= '0';
      ELSIF enb = '1' THEN
        Delay13_out1 <= Delay22_out1;
      END IF;
    END IF;
  END PROCESS Delay13_process;


  Logical_Operator_out1_4 <= Compare_To_Constant1_out1_1 OR Delay13_out1;

  
  Compare_To_Constant_out1_2 <= '1' WHEN Delay18_out1 < to_signed(-16#07F#, 10) ELSE
      '0';

  Constant1_out1_5 <= to_unsigned(16#7F#, 8);

  Delay2_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_2 <= to_unsigned(0, 49);
      ELSIF enb = '1' THEN
        Delay2_out1_2 <= Bit_Concat_out1_1;
      END IF;
    END IF;
  END PROCESS Delay2_2_process;


  
  Compare_To_Zero_out1_1 <= '1' WHEN Delay1_out1_1 < to_signed(16#00#, 6) ELSE
      '0';

  Bit_Slice_out1_1 <= unsigned(Delay1_out1_1(4 DOWNTO 0));

  Shift_Arithmetic_out1 <= Delay2_out1_2 sll to_integer(Bit_Slice_out1_1);

  Bit_Shift_out1 <= SHIFT_RIGHT(Bit_Concat_out1_1, 1);

  Delay3_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1_3 <= to_unsigned(0, 49);
      ELSIF enb = '1' THEN
        Delay3_out1_3 <= Bit_Shift_out1;
      END IF;
    END IF;
  END PROCESS Delay3_3_process;


  
  Switch_out1_5 <= Shift_Arithmetic_out1 WHEN Compare_To_Zero_out1_1 = '0' ELSE
      Delay3_out1_3;

  -- handling denormalized signals
  Constant_out1_2 <= to_signed(-16#07E#, 9);

  Subtract_sub_temp <= resize(Add_out1_1, 32) - resize(Constant_out1_2, 32);
  Subtract_out1_1 <= Subtract_sub_temp(15 DOWNTO 0);

  
  Compare_To_Constant_out1_3 <= '1' WHEN Subtract_out1_1 < to_signed(-16#001F#, 16) ELSE
      '0';

  Subtract_out1_dtc <= Subtract_out1_1(5 DOWNTO 0);

  
  Compare_To_Constant1_out1_2 <= '1' WHEN Subtract_out1_1 > to_signed(16#001F#, 16) ELSE
      '0';

  Constant1_out1_6 <= to_signed(-16#1F#, 6);

  
  Switch_out1_6 <= Subtract_out1_dtc WHEN Compare_To_Constant_out1_3 = '0' ELSE
      Constant1_out1_6;

  Constant2_out1_3 <= to_signed(16#1F#, 6);

  
  Switch1_out1_5 <= Switch_out1_6 WHEN Compare_To_Constant1_out1_2 = '0' ELSE
      Constant2_out1_3;

  Unary_Minus_in0 <=  - (resize(Switch1_out1_5, 7));
  Unary_Minus_out1 <= Unary_Minus_in0(5 DOWNTO 0);

  
  shift_arithmetic_shift_direction <= '1' WHEN Unary_Minus_out1 < to_signed(16#00#, 6) ELSE
      '0';

  Constant_out1_3 <= to_unsigned(16#00000000#, 31);

  Bit_Concat_out1_3 <= Switch_out1_5 & Constant_out1_3;

  
  shift_arithmetic_abs_y <=  - (resize(Unary_Minus_out1, 7)) WHEN Unary_Minus_out1 < to_signed(16#00#, 6) ELSE
      resize(Unary_Minus_out1, 7);
  shift_arithmetic_shift_value <= unsigned(shift_arithmetic_abs_y);

  shift_arithmetic_right <= SHIFT_RIGHT(Bit_Concat_out1_3, to_integer(shift_arithmetic_shift_value));

  shift_arithmetic_left <= Bit_Concat_out1_3 sll to_integer(shift_arithmetic_shift_value);

  
  Shift_Arithmetic_out1_1 <= shift_arithmetic_right WHEN shift_arithmetic_shift_direction = '0' ELSE
      shift_arithmetic_left;

  Bit_Slice1_out1_1 <= Shift_Arithmetic_out1_1(30 DOWNTO 0);

  Bit_Slice_out1_2 <= Shift_Arithmetic_out1_1(79 DOWNTO 31);

  Bit_Set_out1 <= Bit_Slice_out1_2 OR to_unsigned(1, 49);

  
  Switch2_out1_3 <= Bit_Slice_out1_2 WHEN Bit_Slice1_out1_1 = to_unsigned(0, 49) ELSE
      Bit_Set_out1;

  
  Switch1_out1_6 <= Switch_out1_5 WHEN Compare_To_Constant_out1_1 = '0' ELSE
      Switch2_out1_3;

  Bit_Slice_out1_3 <= Switch1_out1_6(47 DOWNTO 0);

  Bit_Slice2_out1_1 <= Bit_Slice_out1_3(23 DOWNTO 22);

  Bit_Slice4_out1_1 <= Bit_Slice2_out1_1(0);

  Bit_Slice1_out1_2 <= Bit_Slice_out1_3(21 DOWNTO 0);

  Bit_Reduce_out1 <= (Bit_Slice1_out1_2(21) OR Bit_Slice1_out1_2(20) OR Bit_Slice1_out1_2(19) OR 
    Bit_Slice1_out1_2(18) OR Bit_Slice1_out1_2(17) OR Bit_Slice1_out1_2(16) OR Bit_Slice1_out1_2(15) OR 
    Bit_Slice1_out1_2(14) OR Bit_Slice1_out1_2(13) OR Bit_Slice1_out1_2(12) OR Bit_Slice1_out1_2(11) OR 
    Bit_Slice1_out1_2(10) OR Bit_Slice1_out1_2(9) OR Bit_Slice1_out1_2(8) OR Bit_Slice1_out1_2(7) OR 
    Bit_Slice1_out1_2(6) OR Bit_Slice1_out1_2(5) OR Bit_Slice1_out1_2(4) OR Bit_Slice1_out1_2(3) OR 
    Bit_Slice1_out1_2(2) OR Bit_Slice1_out1_2(1) OR Bit_Slice1_out1_2(0));

  Bit_Slice5_out1_1 <= Bit_Slice2_out1_1(1);

  Bit_Slice3_out1_1 <= Bit_Slice_out1_3(24);

  Logical_Operator1_out1_3 <= Bit_Slice3_out1_1 OR (Bit_Slice4_out1_1 OR Bit_Reduce_out1);

  Logical_Operator_out1_5 <= Bit_Slice5_out1_1 AND Logical_Operator1_out1_3;

  Delay1_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_2 <= '0';
      ELSIF enb = '1' THEN
        Delay1_out1_2 <= Logical_Operator_out1_5;
      END IF;
    END IF;
  END PROCESS Delay1_2_process;


  Bit_Slice1_out1_3 <= Bit_Slice_out1_3(46 DOWNTO 24);

  reduced_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Bit_Slice1_out1_4 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Bit_Slice1_out1_4 <= Bit_Slice1_out1_3;
      END IF;
    END IF;
  END PROCESS reduced_process;


  Bit_Slice1_out1_dtc <= resize(Bit_Slice1_out1_4, 24);

  Constant_out1_4 <= '1';

  Add_add_cast_1 <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & 
    '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & 
    Constant_out1_4;
  Add_out1_2 <= resize(resize(Bit_Slice1_out1_4, 32) + Add_add_cast_1, 24);

  
  Switch_out1_7 <= Bit_Slice1_out1_dtc WHEN Delay1_out1_2 = '0' ELSE
      Add_out1_2;

  Bit_Slice2_out1_2 <= Switch_out1_7(23);

  Add1_add_cast <= '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & 
    '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & 
    Bit_Slice2_out1_2;
  Add1_out1_1 <= resize(resize(Constant1_out1_5, 32) + Add1_add_cast, 8);

  Add_add_cast_2 <= signed(resize(Add1_out1_1, 32));
  Add_add_temp <= Add_add_cast_2 + resize(Delay18_out1, 32);
  Add_out1_3 <= unsigned(Add_add_temp(7 DOWNTO 0));

  Constant1_out1_7 <= to_unsigned(16#00#, 8);

  
  Switch1_out1_7 <= Add_out1_3 WHEN Compare_To_Constant_out1_2 = '0' ELSE
      Constant1_out1_7;

  Constant4_out1_3 <= to_unsigned(16#FF#, 8);

  
  Switch4_out1_1 <= Switch1_out1_7 WHEN Logical_Operator_out1_4 = '0' ELSE
      Constant4_out1_3;

  
  Switch6_out1_1 <= Constant6_out1 WHEN Relational_Operator_relop1 = '0' ELSE
      Switch4_out1_1;

  Delay1_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay1_out1_3 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay1_out1_3 <= Switch6_out1_1;
      END IF;
    END IF;
  END PROCESS Delay1_3_process;


  Bit_Slice4_out1_2 <= Switch_out1_7(22 DOWNTO 0);

  Bit_Shift_out1_1 <= Bit_Slice4_out1_2 srl 1;

  
  Switch1_out1_8 <= Bit_Slice4_out1_2 WHEN Bit_Slice2_out1_2 = '0' ELSE
      Bit_Shift_out1_1;

  Constant2_out1_4 <= to_unsigned(16#000000#, 23);

  
  Switch2_out1_4 <= Switch1_out1_8 WHEN Compare_To_Constant_out1_2 = '0' ELSE
      Constant2_out1_4;

  Constant5_out1_2 <= to_unsigned(16#000000#, 23);

  Bit_Set_out1_1 <= Switch2_out1_4 OR to_unsigned(16#400000#, 23);

  
  Switch7_out1_1 <= Constant5_out1_2 WHEN Delay13_out1 = '0' ELSE
      Bit_Set_out1_1;

  
  Switch5_out1_1 <= Switch2_out1_4 WHEN Logical_Operator_out1_4 = '0' ELSE
      Switch7_out1_1;

  Delay2_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1_3 <= to_unsigned(16#000000#, 23);
      ELSIF enb = '1' THEN
        Delay2_out1_3 <= Switch5_out1_1;
      END IF;
    END IF;
  END PROCESS Delay2_3_process;


  -- Combine FP sign, exponent, mantissa into 32 bit word
  nfp_out_pack <= Delay_out1 & Delay1_out1_3 & Delay2_out1_3;

  nfp_out <= std_logic_vector(nfp_out_pack);

END rtl;

