LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY my_inverse IS
  PORT( clk                               :   IN    std_logic;
        reset_x                           :   IN    std_logic;
        clk_enable                        :   IN    std_logic;
        en                                :   IN    std_logic;
        in_ri_re                          :   IN    std_logic_vector(31 DOWNTO 0);
        in_ri_im                          :   IN    std_logic_vector(31 DOWNTO 0);
        ce_out                            :   OUT   std_logic;
        valid_out                         :   OUT   std_logic;
        out_ir_re                         :   OUT   std_logic_vector(31 DOWNTO 0);
        out_ir_im                         :   OUT   std_logic_vector(31 DOWNTO 0)
        );
END my_inverse;


ARCHITECTURE rtl OF my_inverse IS

  -- Component Declarations
  COMPONENT func1
    PORT( clk                             :   IN    std_logic;
          reset_x                         :   IN    std_logic;
          enb                             :   IN    std_logic;
          enb_1_1_1                       :   IN    std_logic;
          in1_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          in1_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          in2_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          in2_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          out_re                          :   OUT   std_logic_vector(31 DOWNTO 0);
          out_im                          :   OUT   std_logic_vector(31 DOWNTO 0)
          );
  END COMPONENT;

  COMPONENT func2
    PORT( clk                             :   IN    std_logic;
          reset_x                         :   IN    std_logic;
          enb                             :   IN    std_logic;
          enb_1_1_1                       :   IN    std_logic;
          In1_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          In1_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          In2_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          In2_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          In3_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          In3_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          out_re                          :   OUT   std_logic_vector(31 DOWNTO 0);
          out_im                          :   OUT   std_logic_vector(31 DOWNTO 0)
          );
  END COMPONENT;

  COMPONENT memory
    PORT( clk                             :   IN    std_logic;
          reset_x                         :   IN    std_logic;
          enb                             :   IN    std_logic;
          enb_1_1_1                       :   IN    std_logic;
          din_re                          :   IN    std_logic_vector(31 DOWNTO 0);
          din_im                          :   IN    std_logic_vector(31 DOWNTO 0);
          wr                              :   IN    std_logic;
          add1                            :   IN    std_logic_vector(15 DOWNTO 0);
          add2                            :   IN    std_logic_vector(15 DOWNTO 0);
          add3                            :   IN    std_logic_vector(15 DOWNTO 0);
          out1_re                         :   OUT   std_logic_vector(31 DOWNTO 0);
          out1_im                         :   OUT   std_logic_vector(31 DOWNTO 0);
          out2_re                         :   OUT   std_logic_vector(31 DOWNTO 0);
          out2_im                         :   OUT   std_logic_vector(31 DOWNTO 0);
          out3_re                         :   OUT   std_logic_vector(31 DOWNTO 0);
          out3_im                         :   OUT   std_logic_vector(31 DOWNTO 0)
          );
  END COMPONENT;

  -- Signals
  SIGNAL enb                              : std_logic;
  SIGNAL sit                              : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out          : std_logic;
  SIGNAL intdelay_ctrl_delay_out          : std_logic;
  SIGNAL intdelay_Initial_Val_out         : unsigned(7 DOWNTO 0);
  SIGNAL i_i                              : unsigned(7 DOWNTO 0);
  SIGNAL const_expression                 : unsigned(7 DOWNTO 0);
  SIGNAL i_i_1                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_2                            : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_1               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_2               : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out_1        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_1        : std_logic;
  SIGNAL intdelay_Initial_Val_out_1       : unsigned(7 DOWNTO 0);
  SIGNAL j_j                              : unsigned(7 DOWNTO 0);
  SIGNAL j_j_1                            : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_3               : unsigned(7 DOWNTO 0);
  SIGNAL j_j_2                            : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_4               : unsigned(7 DOWNTO 0);
  SIGNAL sit_1                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_2                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_3                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_4                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_5                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_6                            : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out_2        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_2        : std_logic;
  SIGNAL intdelay_Initial_Val_out_2       : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_5               : unsigned(7 DOWNTO 0);
  SIGNAL k_k                              : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_6               : unsigned(7 DOWNTO 0);
  SIGNAL k_k_1                            : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_7               : unsigned(7 DOWNTO 0);
  SIGNAL k_k_2                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_7                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_8                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_9                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_10                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_11                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_12                           : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_8               : unsigned(7 DOWNTO 0);
  SIGNAL wait_rsvd                        : unsigned(7 DOWNTO 0);
  SIGNAL sit_13                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_14                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_15                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_16                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_17                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_18                           : unsigned(7 DOWNTO 0);
  SIGNAL Unit_Delay2_out1                 : std_logic;
  SIGNAL out0                             : std_logic;
  SIGNAL intdelay_ctrl_const_out_3        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_3        : std_logic;
  SIGNAL intdelay_Initial_Val_out_3       : unsigned(7 DOWNTO 0);
  SIGNAL i1                               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_9               : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out_4        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_4        : std_logic;
  SIGNAL intdelay_Initial_Val_out_4       : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_10              : unsigned(7 DOWNTO 0);
  SIGNAL sit_19                           : unsigned(7 DOWNTO 0);
  SIGNAL j1                               : unsigned(7 DOWNTO 0);
  SIGNAL j1_1                             : unsigned(7 DOWNTO 0);
  SIGNAL j1_2                             : unsigned(7 DOWNTO 0);
  SIGNAL j1_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_1                           : std_logic;
  SIGNAL out0_2                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_3                           : std_logic;
  SIGNAL out0_4                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_5                           : std_logic;
  SIGNAL out0_6                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_7                           : std_logic;
  SIGNAL out0_8                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_9                           : std_logic;
  SIGNAL out0_10                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_11                          : std_logic;
  SIGNAL out0_12                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_13                          : std_logic;
  SIGNAL out0_14                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_15                          : std_logic;
  SIGNAL out0_16                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_17                          : std_logic;
  SIGNAL out0_18                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_19                          : std_logic;
  SIGNAL out0_20                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_21                          : std_logic;
  SIGNAL out0_22                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_23                          : std_logic;
  SIGNAL out0_24                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_25                          : std_logic;
  SIGNAL out0_26                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_27                          : std_logic;
  SIGNAL out0_28                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_29                          : std_logic;
  SIGNAL out0_30                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_31                          : std_logic;
  SIGNAL j1_4                             : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out                     : unsigned(7 DOWNTO 0);
  SIGNAL out0_32                          : std_logic;
  SIGNAL i1_1                             : unsigned(7 DOWNTO 0);
  SIGNAL i1_2                             : unsigned(7 DOWNTO 0);
  SIGNAL i1_3                             : unsigned(7 DOWNTO 0);
  SIGNAL i1_4                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_33                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_34                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_35                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_36                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_37                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_38                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_39                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_40                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_41                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_42                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_43                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_44                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_45                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_46                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_47                          : unsigned(7 DOWNTO 0);
  SIGNAL i1_5                             : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out_1                   : unsigned(7 DOWNTO 0);
  SIGNAL out0_48                          : std_logic;
  SIGNAL sit_20                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_21                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_22                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_49                          : std_logic;
  SIGNAL sit_23                           : unsigned(7 DOWNTO 0);
  SIGNAL wait_rsvd_1                      : unsigned(7 DOWNTO 0);
  SIGNAL wait_rsvd_2                      : unsigned(7 DOWNTO 0);
  SIGNAL out0_50                          : std_logic;
  SIGNAL wait_rsvd_3                      : unsigned(7 DOWNTO 0);
  SIGNAL out0_51                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_52                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_53                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_54                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_55                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_56                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_57                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_58                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_59                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_60                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_61                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_62                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_63                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_64                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_65                          : unsigned(7 DOWNTO 0);
  SIGNAL wait_rsvd_4                      : unsigned(7 DOWNTO 0);
  SIGNAL sit_24                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_66                          : std_logic;
  SIGNAL sit_25                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_67                          : std_logic;
  SIGNAL sit_26                           : unsigned(7 DOWNTO 0);
  SIGNAL k_k_3                            : unsigned(7 DOWNTO 0);
  SIGNAL k_k_4                            : unsigned(7 DOWNTO 0);
  SIGNAL k_k_5                            : unsigned(7 DOWNTO 0);
  SIGNAL k_k_6                            : unsigned(7 DOWNTO 0);
  SIGNAL k_k_7                            : unsigned(7 DOWNTO 0);
  SIGNAL k_k_8                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_68                          : std_logic;
  SIGNAL k_k_9                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_69                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_70                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_71                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_72                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_73                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_74                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_75                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_76                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_77                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_78                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_79                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_80                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_81                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_82                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_83                          : unsigned(7 DOWNTO 0);
  SIGNAL k_k_10                           : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out_2                   : unsigned(7 DOWNTO 0);
  SIGNAL sit_27                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_84                          : std_logic;
  SIGNAL sit_28                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_85                          : std_logic;
  SIGNAL sit_29                           : unsigned(7 DOWNTO 0);
  SIGNAL j_j_3                            : unsigned(7 DOWNTO 0);
  SIGNAL j_j_4                            : unsigned(7 DOWNTO 0);
  SIGNAL j_j_5                            : unsigned(7 DOWNTO 0);
  SIGNAL j_j_6                            : unsigned(7 DOWNTO 0);
  SIGNAL j_j_7                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_86                          : std_logic;
  SIGNAL j_j_8                            : unsigned(7 DOWNTO 0);
  SIGNAL j_j_9                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_87                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_88                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_89                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_90                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_91                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_92                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_93                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_94                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_95                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_96                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_97                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_98                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_99                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_100                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_101                         : unsigned(7 DOWNTO 0);
  SIGNAL j_j_10                           : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out_3                   : unsigned(7 DOWNTO 0);
  SIGNAL i_i_3                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_4                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_5                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_6                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_7                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_102                         : std_logic;
  SIGNAL i_i_8                            : unsigned(7 DOWNTO 0);
  SIGNAL i_i_9                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_103                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_104                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_105                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_106                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_107                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_108                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_109                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_110                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_111                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_112                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_113                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_114                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_115                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_116                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_117                         : unsigned(7 DOWNTO 0);
  SIGNAL i_i_10                           : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out_4                   : unsigned(7 DOWNTO 0);
  SIGNAL sit_30                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_118                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_119                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_120                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_121                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_122                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_123                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_124                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_125                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_126                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_127                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_128                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_129                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_130                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_131                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_132                         : unsigned(7 DOWNTO 0);
  SIGNAL sit_out                          : unsigned(7 DOWNTO 0);
  SIGNAL valid_out_1                      : std_logic;
  SIGNAL valid_out_2                      : std_logic;
  SIGNAL out0_133                         : std_logic;
  SIGNAL valid_out_3                      : std_logic;
  SIGNAL out0_134                         : std_logic;
  SIGNAL valid_out_4                      : std_logic;
  SIGNAL out0_135                         : std_logic;
  SIGNAL valid_out_5                      : std_logic;
  SIGNAL out0_136                         : std_logic;
  SIGNAL valid_out_6                      : std_logic;
  SIGNAL out0_137                         : std_logic;
  SIGNAL valid_out_7                      : std_logic;
  SIGNAL out0_138                         : std_logic;
  SIGNAL valid_out_8                      : std_logic;
  SIGNAL out0_139                         : std_logic;
  SIGNAL valid_out_9                      : std_logic;
  SIGNAL out0_140                         : std_logic;
  SIGNAL valid_out_10                     : std_logic;
  SIGNAL out0_141                         : std_logic;
  SIGNAL valid_out_11                     : std_logic;
  SIGNAL out0_142                         : std_logic;
  SIGNAL valid_out_12                     : std_logic;
  SIGNAL out0_143                         : std_logic;
  SIGNAL valid_out_13                     : std_logic;
  SIGNAL out0_144                         : std_logic;
  SIGNAL valid_out_14                     : std_logic;
  SIGNAL out0_145                         : std_logic;
  SIGNAL valid_out_15                     : std_logic;
  SIGNAL out0_146                         : std_logic;
  SIGNAL valid_out_16                     : std_logic;
  SIGNAL out0_147                         : std_logic;
  SIGNAL valid_out_17                     : std_logic;
  SIGNAL valid_out_18                     : std_logic;
  SIGNAL Unit_Delay4_out1                 : std_logic;
  SIGNAL Data_Type_Conversion_out1        : std_logic;
  SIGNAL data_out_re                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_1                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_1                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_2                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_2                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_1                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_1                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_3                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_3                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_2                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_2                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_4                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_4                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_3                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_3                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL relop1_relop1                    : std_logic;
  SIGNAL ram_out_re_5                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_5                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL relop_relop1                     : std_logic;
  SIGNAL ram_out_re_6                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_6                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_7                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_7                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_8                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_8                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_9                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_9                     : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_10                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_10                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_11                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_11                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_12                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_12                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_13                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_13                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_14                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_14                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_15                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_15                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL Unit_Delay3_out1_re              : std_logic_vector(31 DOWNTO 0);
  SIGNAL Unit_Delay3_out1_im              : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_16                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_16                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL we                               : std_logic;
  SIGNAL we_1                             : std_logic;
  SIGNAL out0_148                         : std_logic;
  SIGNAL we_2                             : std_logic;
  SIGNAL out0_149                         : std_logic;
  SIGNAL we_3                             : std_logic;
  SIGNAL out0_150                         : std_logic;
  SIGNAL we_4                             : std_logic;
  SIGNAL out0_151                         : std_logic;
  SIGNAL we_5                             : std_logic;
  SIGNAL we_6                             : std_logic;
  SIGNAL we_7                             : std_logic;
  SIGNAL out0_152                         : std_logic;
  SIGNAL we_8                             : std_logic;
  SIGNAL out0_153                         : std_logic;
  SIGNAL we_9                             : std_logic;
  SIGNAL out0_154                         : std_logic;
  SIGNAL we_10                            : std_logic;
  SIGNAL out0_155                         : std_logic;
  SIGNAL we_11                            : std_logic;
  SIGNAL out0_156                         : std_logic;
  SIGNAL we_12                            : std_logic;
  SIGNAL out0_157                         : std_logic;
  SIGNAL we_13                            : std_logic;
  SIGNAL out0_158                         : std_logic;
  SIGNAL we_14                            : std_logic;
  SIGNAL out0_159                         : std_logic;
  SIGNAL we_15                            : std_logic;
  SIGNAL out0_160                         : std_logic;
  SIGNAL we_16                            : std_logic;
  SIGNAL out0_161                         : std_logic;
  SIGNAL we_17                            : std_logic;
  SIGNAL out0_162                         : std_logic;
  SIGNAL we_18                            : std_logic;
  SIGNAL we_19                            : std_logic;
  SIGNAL we_20                            : std_logic;
  SIGNAL we_21                            : std_logic;
  SIGNAL ram_add1                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_11                           : unsigned(15 DOWNTO 0);
  SIGNAL jj                               : unsigned(15 DOWNTO 0);
  SIGNAL i_i_11                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_1                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_163                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_12                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_1                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_12                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_2                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_164                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_3                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_165                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_4                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_166                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_5                       : unsigned(15 DOWNTO 0);
  SIGNAL j_j_13                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_2                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_13                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_6                       : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_7                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_167                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_14                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_3                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_14                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_8                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_168                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_15                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_4                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_15                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_9                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_169                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_10                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_170                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_16                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_5                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_16                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_11                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_171                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_12                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_172                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_13                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_173                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_17                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_6                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_17                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_14                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_174                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_15                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_175                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_18                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_7                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_18                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_16                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_176                         : unsigned(15 DOWNTO 0);
  SIGNAL n_n                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_177                         : unsigned(7 DOWNTO 0);
  SIGNAL j_j_19                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_8                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_19                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_17                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_178                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_18                      : unsigned(15 DOWNTO 0);
  SIGNAL j_j_20                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_9                             : unsigned(15 DOWNTO 0);
  SIGNAL i_i_20                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_19                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_20                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add1_21                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_21                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_10                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_21                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_1                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_179                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_22                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_11                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_22                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_2                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_180                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_3                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_181                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_4                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_182                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_5                       : unsigned(15 DOWNTO 0);
  SIGNAL j_j_23                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_12                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_23                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_6                       : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_7                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_183                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_24                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_13                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_24                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_8                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_184                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_25                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_14                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_25                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_9                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_185                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_10                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_186                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_26                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_15                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_26                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_11                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_187                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_12                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_188                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_13                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_189                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_27                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_16                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_27                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_14                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_190                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_15                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_191                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_28                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_17                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_28                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_16                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_192                         : unsigned(15 DOWNTO 0);
  SIGNAL n_n_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_193                         : unsigned(7 DOWNTO 0);
  SIGNAL j_j_29                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_18                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_29                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_17                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_194                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_18                      : unsigned(15 DOWNTO 0);
  SIGNAL j_j_30                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_19                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_30                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_19                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_20                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add2_21                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_31                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_20                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_31                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_1                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_195                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_32                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_21                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_32                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_2                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_196                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_3                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_197                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_4                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_198                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_5                       : unsigned(15 DOWNTO 0);
  SIGNAL j_j_33                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_22                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_33                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_6                       : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_7                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_199                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_34                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_23                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_34                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_8                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_200                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_35                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_24                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_35                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_9                       : unsigned(15 DOWNTO 0);
  SIGNAL out0_201                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_10                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_202                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_36                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_25                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_36                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_11                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_203                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_12                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_204                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_13                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_205                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_37                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_26                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_37                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_14                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_206                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_15                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_207                         : unsigned(15 DOWNTO 0);
  SIGNAL j_j_38                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_27                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_38                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_16                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_208                         : unsigned(15 DOWNTO 0);
  SIGNAL n_n_2                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_209                         : unsigned(7 DOWNTO 0);
  SIGNAL j_j_39                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_28                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_39                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_17                      : unsigned(15 DOWNTO 0);
  SIGNAL out0_210                         : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_18                      : unsigned(15 DOWNTO 0);
  SIGNAL j_j_40                           : unsigned(15 DOWNTO 0);
  SIGNAL jj_29                            : unsigned(15 DOWNTO 0);
  SIGNAL i_i_40                           : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_19                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_20                      : unsigned(15 DOWNTO 0);
  SIGNAL ram_add3_21                      : unsigned(15 DOWNTO 0);
  SIGNAL dout2_re                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout2_im                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL p2_re                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p2_im                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_4                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_4                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_5                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_5                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_6                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_6                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_7                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_7                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_8                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_8                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_9                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_9                        : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_10                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_10                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_11                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_11                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_12                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_12                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_13                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_13                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out1_re                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out1_im                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_14                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_14                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_15                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_15                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_16                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_16                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_17                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_17                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_18                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_18                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout1_re                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout1_im                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL p1_re                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p1_im                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_19                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_19                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_20                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_20                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_21                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_21                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_22                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_22                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_23                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_23                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_24                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_24                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_25                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_25                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_26                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_26                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_27                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_27                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_28                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_28                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_29                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_29                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_30                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_30                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_31                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_31                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_32                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_32                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_33                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_33                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL func1_out1_re                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL func1_out1_im                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL p5_re                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p5_im                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out3_re                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out3_im                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL p5_re_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL p5_im_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout5_re                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout5_im                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_34                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_34                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_35                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_35                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_36                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_36                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_37                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_37                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_38                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_38                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_39                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_39                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_40                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_40                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_41                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_41                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_42                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_42                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_43                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_43                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_44                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_44                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_45                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_45                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_46                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_46                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_47                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_47                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_48                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_48                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL p4_re                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p4_im                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out2_re                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL memory_out2_im                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL p4_re_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL p4_im_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout4_re                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout4_im                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_49                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_49                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_50                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_50                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_51                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_51                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_52                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_52                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_53                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_53                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_54                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_54                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_55                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_55                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_56                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_56                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_57                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_57                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_58                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_58                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_59                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_59                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_60                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_60                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_61                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_61                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_62                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_62                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_63                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_63                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL p3_re                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p3_im                            : std_logic_vector(31 DOWNTO 0);
  SIGNAL p3_re_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL p3_im_1                          : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout3_re                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL dout3_im                         : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_64                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_64                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_65                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_65                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_66                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_66                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_67                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_67                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_68                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_68                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_69                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_69                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_70                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_70                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_71                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_71                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_72                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_72                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_73                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_73                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_74                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_74                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_75                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_75                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_76                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_76                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_77                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_77                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_78                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_78                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL func2_out1_re                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL func2_out1_im                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_17                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_17                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_79                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_79                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_80                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_80                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_81                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_81                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_82                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_82                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_83                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_83                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_84                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_84                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_85                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_85                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_86                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_86                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_87                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_87                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_88                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_88                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_89                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_89                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_re_18                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL ram_out_im_18                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_90                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_90                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_1                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_1                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_91                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_91                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_2                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_2                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_92                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_92                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_3                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_3                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_93                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_93                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_4                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_4                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_94                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_94                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_5                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_5                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_95                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_95                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_6                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_6                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_96                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_96                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_7                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_7                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_97                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_97                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_8                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_8                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_98                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_98                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_9                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_9                    : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_99                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_99                       : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_10                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_10                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_100                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_100                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_11                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_11                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_101                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_101                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_12                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_12                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_102                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_102                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_13                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_13                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_103                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_103                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_14                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_14                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_re_104                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL out0_im_104                      : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_15                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_15                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_re_16                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL data_out_im_16                   : std_logic_vector(31 DOWNTO 0);
  SIGNAL Unit_Delay1_out1_re              : std_logic_vector(31 DOWNTO 0);
  SIGNAL Unit_Delay1_out1_im              : std_logic_vector(31 DOWNTO 0);

BEGIN
  Ufunc1_1 : func1
    PORT MAP( clk => clk,
              reset_x => reset_x,
              enb => clk_enable,
              enb_1_1_1 => clk_enable,
              in1_re => dout1_re,
              in1_im => dout1_im,
              in2_re => dout2_re,
              in2_im => dout2_im,
              out_re => func1_out1_re,
              out_im => func1_out1_im
              );

  Ufunc2_1 : func2
    PORT MAP( clk => clk,
              reset_x => reset_x,
              enb => clk_enable,
              enb_1_1_1 => clk_enable,
              In1_re => dout3_re,
              In1_im => dout3_im,
              In2_re => dout4_re,
              In2_im => dout4_im,
              In3_re => dout5_re,
              In3_im => dout5_im,
              out_re => func2_out1_re,
              out_im => func2_out1_im
              );

  Umemory_1 : memory
    PORT MAP( clk => clk,
              reset_x => reset_x,
              enb => clk_enable,
              enb_1_1_1 => clk_enable,
              din_re => ram_out_re_18,
              din_im => ram_out_im_18,
              wr => we_21,
              add1 => std_logic_vector(ram_add1_21),
              add2 => std_logic_vector(ram_add2_21),
              add3 => std_logic_vector(ram_add3_21),
              out1_re => memory_out1_re,
              out1_im => memory_out1_im,
              out2_re => memory_out2_re,
              out2_im => memory_out2_im,
              out3_re => memory_out3_re,
              out3_im => memory_out3_im
              );

  sit <= to_unsigned(16#00#, 8);

  intdelay_ctrl_const_out <= '1';

  enb <= clk_enable;

  intdelay_ctrl_delay_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out <= intdelay_ctrl_const_out;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay_process;


  intdelay_Initial_Val_out <= to_unsigned(16#01#, 8);

  i_i <= to_unsigned(16#01#, 8);

  const_expression <= to_unsigned(16#01#, 8);

  i_i_1 <= to_unsigned(16#01#, 8);

  i_i_2 <= to_unsigned(16#01#, 8);

  const_expression_1 <= to_unsigned(16#01#, 8);

  const_expression_2 <= to_unsigned(16#01#, 8);

  intdelay_ctrl_const_out_1 <= '1';

  intdelay_ctrl_delay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_1 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_1 <= intdelay_ctrl_const_out_1;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay1_process;


  intdelay_Initial_Val_out_1 <= to_unsigned(16#01#, 8);

  j_j <= to_unsigned(16#11#, 8);

  j_j_1 <= to_unsigned(16#11#, 8);

  const_expression_3 <= to_unsigned(16#01#, 8);

  j_j_2 <= to_unsigned(16#01#, 8);

  const_expression_4 <= to_unsigned(16#01#, 8);

  sit_1 <= to_unsigned(16#00#, 8);

  sit_2 <= to_unsigned(16#0C#, 8);

  sit_3 <= to_unsigned(16#02#, 8);

  sit_4 <= to_unsigned(16#0B#, 8);

  sit_5 <= to_unsigned(16#05#, 8);

  sit_6 <= to_unsigned(16#0A#, 8);

  intdelay_ctrl_const_out_2 <= '1';

  intdelay_ctrl_delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_2 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_2 <= intdelay_ctrl_const_out_2;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay2_process;


  intdelay_Initial_Val_out_2 <= to_unsigned(16#01#, 8);

  const_expression_5 <= to_unsigned(16#01#, 8);

  k_k <= to_unsigned(16#01#, 8);

  const_expression_6 <= to_unsigned(16#01#, 8);

  k_k_1 <= to_unsigned(16#01#, 8);

  const_expression_7 <= to_unsigned(16#01#, 8);

  k_k_2 <= to_unsigned(16#01#, 8);

  sit_7 <= to_unsigned(16#09#, 8);

  sit_8 <= to_unsigned(16#08#, 8);

  sit_9 <= to_unsigned(16#06#, 8);

  sit_10 <= to_unsigned(16#03#, 8);

  sit_11 <= to_unsigned(16#05#, 8);

  sit_12 <= to_unsigned(16#04#, 8);

  const_expression_8 <= to_unsigned(16#01#, 8);

  wait_rsvd <= to_unsigned(16#00#, 8);

  sit_13 <= to_unsigned(16#27#, 8);

  sit_14 <= to_unsigned(16#20#, 8);

  sit_15 <= to_unsigned(16#1F#, 8);

  sit_16 <= to_unsigned(16#03#, 8);

  sit_17 <= to_unsigned(16#15#, 8);

  sit_18 <= to_unsigned(16#02#, 8);

  Unit_Delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Unit_Delay2_out1 <= '0';
      ELSIF enb = '1' THEN
        Unit_Delay2_out1 <= en;
      END IF;
    END IF;
  END PROCESS Unit_Delay2_process;


  
  out0 <= '1' WHEN Unit_Delay2_out1 = '1' ELSE
      '0';

  intdelay_ctrl_const_out_3 <= '1';

  intdelay_ctrl_delay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_3 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_3 <= intdelay_ctrl_const_out_3;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay3_process;


  intdelay_Initial_Val_out_3 <= to_unsigned(16#01#, 8);

  i1 <= to_unsigned(16#01#, 8);

  const_expression_9 <= to_unsigned(16#01#, 8);

  intdelay_ctrl_const_out_4 <= '1';

  intdelay_ctrl_delay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_4 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_4 <= intdelay_ctrl_const_out_4;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay4_process;


  intdelay_Initial_Val_out_4 <= to_unsigned(16#01#, 8);

  const_expression_10 <= to_unsigned(16#01#, 8);

  sit_19 <= to_unsigned(16#01#, 8);

  j1_1 <= j1 + const_expression_10;

  
  j1_3 <= j1 WHEN out0 = '0' ELSE
      j1_2;

  
  out0_2 <= j1 WHEN out0_1 = '0' ELSE
      j1;

  
  out0_4 <= out0_2 WHEN out0_3 = '0' ELSE
      j1;

  
  out0_6 <= out0_4 WHEN out0_5 = '0' ELSE
      j1;

  
  out0_8 <= out0_6 WHEN out0_7 = '0' ELSE
      j1;

  
  out0_10 <= out0_8 WHEN out0_9 = '0' ELSE
      j1;

  
  out0_12 <= out0_10 WHEN out0_11 = '0' ELSE
      j1;

  
  out0_14 <= out0_12 WHEN out0_13 = '0' ELSE
      j1;

  
  out0_16 <= out0_14 WHEN out0_15 = '0' ELSE
      j1;

  
  out0_18 <= out0_16 WHEN out0_17 = '0' ELSE
      j1;

  
  out0_20 <= out0_18 WHEN out0_19 = '0' ELSE
      j1;

  
  out0_22 <= out0_20 WHEN out0_21 = '0' ELSE
      j1;

  
  out0_24 <= out0_22 WHEN out0_23 = '0' ELSE
      j1;

  
  out0_26 <= out0_24 WHEN out0_25 = '0' ELSE
      j1;

  
  out0_28 <= out0_26 WHEN out0_27 = '0' ELSE
      j1;

  
  out0_30 <= out0_28 WHEN out0_29 = '0' ELSE
      j1;

  
  j1_4 <= out0_30 WHEN out0_31 = '0' ELSE
      j1_3;

  intdelay5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out <= j1_4;
      END IF;
    END IF;
  END PROCESS intdelay5_process;


  
  j1 <= intdelay_Initial_Val_out_4 WHEN intdelay_ctrl_delay_out_4 = '0' ELSE
      intdelay_out;

  
  i1_2 <= i1_1 WHEN out0_32 = '0' ELSE
      i1;

  
  i1_4 <= i1_3 WHEN out0 = '0' ELSE
      i1_2;

  
  out0_33 <= i1_3 WHEN out0_1 = '0' ELSE
      i1_3;

  
  out0_34 <= out0_33 WHEN out0_3 = '0' ELSE
      i1_3;

  
  out0_35 <= out0_34 WHEN out0_5 = '0' ELSE
      i1_3;

  
  out0_36 <= out0_35 WHEN out0_7 = '0' ELSE
      i1_3;

  
  out0_37 <= out0_36 WHEN out0_9 = '0' ELSE
      i1_3;

  
  out0_38 <= out0_37 WHEN out0_11 = '0' ELSE
      i1_3;

  
  out0_39 <= out0_38 WHEN out0_13 = '0' ELSE
      i1_3;

  
  out0_40 <= out0_39 WHEN out0_15 = '0' ELSE
      i1_3;

  
  out0_41 <= out0_40 WHEN out0_17 = '0' ELSE
      i1_3;

  
  out0_42 <= out0_41 WHEN out0_19 = '0' ELSE
      i1_3;

  
  out0_43 <= out0_42 WHEN out0_21 = '0' ELSE
      i1_3;

  
  out0_44 <= out0_43 WHEN out0_23 = '0' ELSE
      i1_3;

  
  out0_45 <= out0_44 WHEN out0_25 = '0' ELSE
      i1_3;

  
  out0_46 <= out0_45 WHEN out0_27 = '0' ELSE
      i1_3;

  
  out0_47 <= out0_46 WHEN out0_29 = '0' ELSE
      i1_3;

  
  i1_5 <= out0_47 WHEN out0_31 = '0' ELSE
      i1_4;

  intdelay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_1 <= i1_5;
      END IF;
    END IF;
  END PROCESS intdelay4_process;


  
  i1_3 <= intdelay_Initial_Val_out_3 WHEN intdelay_ctrl_delay_out_3 = '0' ELSE
      intdelay_out_1;

  i1_1 <= i1_3 + const_expression_9;

  
  out0_32 <= '1' WHEN i1_1 > to_unsigned(16#10#, 8) ELSE
      '0';

  
  j1_2 <= j1 WHEN out0_32 = '0' ELSE
      j1_1;

  
  out0_48 <= '1' WHEN j1_2 > to_unsigned(16#10#, 8) ELSE
      '0';

  
  sit_21 <= sit_20 WHEN out0_48 = '0' ELSE
      sit_19;

  
  sit_22 <= sit_20 WHEN out0 = '0' ELSE
      sit_21;

  
  sit_23 <= sit_18 WHEN out0_49 = '0' ELSE
      sit_20;

  wait_rsvd_2 <= wait_rsvd_1 + const_expression_8;

  
  wait_rsvd_3 <= wait_rsvd_2 WHEN out0_50 = '0' ELSE
      wait_rsvd;

  
  out0_51 <= wait_rsvd_1 WHEN out0_1 = '0' ELSE
      wait_rsvd_1;

  
  out0_52 <= out0_51 WHEN out0_3 = '0' ELSE
      wait_rsvd_1;

  
  out0_53 <= out0_52 WHEN out0_5 = '0' ELSE
      wait_rsvd_1;

  
  out0_54 <= out0_53 WHEN out0_7 = '0' ELSE
      wait_rsvd_1;

  
  out0_55 <= out0_54 WHEN out0_9 = '0' ELSE
      wait_rsvd_1;

  
  out0_56 <= out0_55 WHEN out0_11 = '0' ELSE
      wait_rsvd_1;

  
  out0_57 <= out0_56 WHEN out0_13 = '0' ELSE
      wait_rsvd_1;

  
  out0_58 <= out0_57 WHEN out0_15 = '0' ELSE
      wait_rsvd_1;

  
  out0_59 <= out0_58 WHEN out0_17 = '0' ELSE
      wait_rsvd_1;

  
  out0_60 <= out0_59 WHEN out0_19 = '0' ELSE
      wait_rsvd_3;

  
  out0_61 <= out0_60 WHEN out0_21 = '0' ELSE
      wait_rsvd_1;

  
  out0_62 <= out0_61 WHEN out0_23 = '0' ELSE
      wait_rsvd_1;

  
  out0_63 <= out0_62 WHEN out0_25 = '0' ELSE
      wait_rsvd_1;

  
  out0_64 <= out0_63 WHEN out0_27 = '0' ELSE
      wait_rsvd_1;

  
  out0_65 <= out0_64 WHEN out0_29 = '0' ELSE
      wait_rsvd_1;

  
  wait_rsvd_4 <= out0_65 WHEN out0_31 = '0' ELSE
      wait_rsvd_1;

  intdelay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        wait_rsvd_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        wait_rsvd_1 <= wait_rsvd_4;
      END IF;
    END IF;
  END PROCESS intdelay2_process;


  
  out0_50 <= '1' WHEN wait_rsvd_1 = to_unsigned(16#11#, 8) ELSE
      '0';

  
  sit_24 <= sit_20 WHEN out0_50 = '0' ELSE
      sit_13;

  
  sit_25 <= sit_10 WHEN out0_66 = '0' ELSE
      sit_11;

  
  sit_26 <= sit_20 WHEN out0_67 = '0' ELSE
      sit_8;

  k_k_4 <= k_k_3 + const_expression_7;

  
  out0_66 <= '1' WHEN k_k_3 = to_unsigned(16#20#, 8) ELSE
      '0';

  
  k_k_5 <= k_k_4 WHEN out0_66 = '0' ELSE
      k_k_2;

  k_k_6 <= k_k_3 + const_expression_6;

  
  out0_67 <= '1' WHEN k_k_3 = to_unsigned(16#20#, 8) ELSE
      '0';

  
  k_k_7 <= k_k_6 WHEN out0_67 = '0' ELSE
      k_k_1;

  k_k_8 <= k_k_3 + const_expression_5;

  
  k_k_9 <= k_k_8 WHEN out0_68 = '0' ELSE
      k_k;

  
  out0_69 <= k_k_3 WHEN out0_1 = '0' ELSE
      k_k_3;

  
  out0_70 <= out0_69 WHEN out0_3 = '0' ELSE
      k_k_3;

  
  out0_71 <= out0_70 WHEN out0_5 = '0' ELSE
      k_k_3;

  
  out0_72 <= out0_71 WHEN out0_7 = '0' ELSE
      k_k_3;

  
  out0_73 <= out0_72 WHEN out0_9 = '0' ELSE
      k_k_9;

  
  out0_74 <= out0_73 WHEN out0_11 = '0' ELSE
      k_k_7;

  
  out0_75 <= out0_74 WHEN out0_13 = '0' ELSE
      k_k_3;

  
  out0_76 <= out0_75 WHEN out0_15 = '0' ELSE
      k_k_5;

  
  out0_77 <= out0_76 WHEN out0_17 = '0' ELSE
      k_k_3;

  
  out0_78 <= out0_77 WHEN out0_19 = '0' ELSE
      k_k_3;

  
  out0_79 <= out0_78 WHEN out0_21 = '0' ELSE
      k_k_3;

  
  out0_80 <= out0_79 WHEN out0_23 = '0' ELSE
      k_k_3;

  
  out0_81 <= out0_80 WHEN out0_25 = '0' ELSE
      k_k_3;

  
  out0_82 <= out0_81 WHEN out0_27 = '0' ELSE
      k_k_3;

  
  out0_83 <= out0_82 WHEN out0_29 = '0' ELSE
      k_k_3;

  
  k_k_10 <= out0_83 WHEN out0_31 = '0' ELSE
      k_k_3;

  intdelay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_2 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_2 <= k_k_10;
      END IF;
    END IF;
  END PROCESS intdelay1_process;


  
  k_k_3 <= intdelay_Initial_Val_out_2 WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2;

  
  out0_68 <= '1' WHEN k_k_3 = to_unsigned(16#20#, 8) ELSE
      '0';

  
  sit_27 <= sit_20 WHEN out0_68 = '0' ELSE
      sit_7;

  
  sit_28 <= sit_5 WHEN out0_84 = '0' ELSE
      sit_6;

  
  sit_29 <= sit_3 WHEN out0_85 = '0' ELSE
      sit_4;

  j_j_4 <= j_j_3 + const_expression_4;

  j_j_5 <= j_j_3 + const_expression_3;

  
  out0_84 <= '1' WHEN j_j_5 > to_unsigned(16#10#, 8) ELSE
      '0';

  
  j_j_6 <= j_j_5 WHEN out0_84 = '0' ELSE
      j_j_2;

  
  j_j_7 <= j_j_3 WHEN out0_85 = '0' ELSE
      j_j_1;

  
  j_j_9 <= j_j_8 WHEN out0_86 = '0' ELSE
      j_j;

  
  out0_87 <= j_j_3 WHEN out0_1 = '0' ELSE
      j_j_9;

  
  out0_88 <= out0_87 WHEN out0_3 = '0' ELSE
      j_j_3;

  
  out0_89 <= out0_88 WHEN out0_5 = '0' ELSE
      j_j_7;

  
  out0_90 <= out0_89 WHEN out0_7 = '0' ELSE
      j_j_6;

  
  out0_91 <= out0_90 WHEN out0_9 = '0' ELSE
      j_j_3;

  
  out0_92 <= out0_91 WHEN out0_11 = '0' ELSE
      j_j_3;

  
  out0_93 <= out0_92 WHEN out0_13 = '0' ELSE
      j_j_3;

  
  out0_94 <= out0_93 WHEN out0_15 = '0' ELSE
      j_j_3;

  
  out0_95 <= out0_94 WHEN out0_17 = '0' ELSE
      j_j_3;

  
  out0_96 <= out0_95 WHEN out0_19 = '0' ELSE
      j_j_3;

  
  out0_97 <= out0_96 WHEN out0_21 = '0' ELSE
      j_j_3;

  
  out0_98 <= out0_97 WHEN out0_23 = '0' ELSE
      j_j_3;

  
  out0_99 <= out0_98 WHEN out0_25 = '0' ELSE
      j_j_3;

  
  out0_100 <= out0_99 WHEN out0_27 = '0' ELSE
      j_j_3;

  
  out0_101 <= out0_100 WHEN out0_29 = '0' ELSE
      j_j_3;

  
  j_j_10 <= out0_101 WHEN out0_31 = '0' ELSE
      j_j_3;

  intdelay_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_3 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_3 <= j_j_10;
      END IF;
    END IF;
  END PROCESS intdelay_process;


  
  j_j_3 <= intdelay_Initial_Val_out_1 WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_3;

  i_i_4 <= i_i_3 + const_expression_1;

  
  out0_49 <= '1' WHEN i_i_3 <= to_unsigned(16#10#, 8) ELSE
      '0';

  
  i_i_5 <= i_i_2 WHEN out0_49 = '0' ELSE
      i_i_4;

  i_i_6 <= i_i_3 + const_expression;

  
  out0_85 <= '1' WHEN i_i_6 > to_unsigned(16#10#, 8) ELSE
      '0';

  
  i_i_7 <= i_i_6 WHEN out0_85 = '0' ELSE
      i_i_1;

  
  i_i_9 <= i_i_8 WHEN out0_102 = '0' ELSE
      i_i;

  
  out0_103 <= i_i_3 WHEN out0_1 = '0' ELSE
      i_i_9;

  
  out0_104 <= out0_103 WHEN out0_3 = '0' ELSE
      i_i_3;

  
  out0_105 <= out0_104 WHEN out0_5 = '0' ELSE
      i_i_7;

  
  out0_106 <= out0_105 WHEN out0_7 = '0' ELSE
      i_i_3;

  
  out0_107 <= out0_106 WHEN out0_9 = '0' ELSE
      i_i_3;

  
  out0_108 <= out0_107 WHEN out0_11 = '0' ELSE
      i_i_3;

  
  out0_109 <= out0_108 WHEN out0_13 = '0' ELSE
      i_i_3;

  
  out0_110 <= out0_109 WHEN out0_15 = '0' ELSE
      i_i_3;

  
  out0_111 <= out0_110 WHEN out0_17 = '0' ELSE
      i_i_3;

  
  out0_112 <= out0_111 WHEN out0_19 = '0' ELSE
      i_i_3;

  
  out0_113 <= out0_112 WHEN out0_21 = '0' ELSE
      i_i_3;

  
  out0_114 <= out0_113 WHEN out0_23 = '0' ELSE
      i_i_3;

  
  out0_115 <= out0_114 WHEN out0_25 = '0' ELSE
      i_i_3;

  
  out0_116 <= out0_115 WHEN out0_27 = '0' ELSE
      i_i_3;

  
  out0_117 <= out0_116 WHEN out0_29 = '0' ELSE
      i_i_5;

  
  i_i_10 <= out0_117 WHEN out0_31 = '0' ELSE
      i_i_3;

  intdelay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_4 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_4 <= i_i_10;
      END IF;
    END IF;
  END PROCESS intdelay3_process;


  
  i_i_3 <= intdelay_Initial_Val_out WHEN intdelay_ctrl_delay_out = '0' ELSE
      intdelay_out_4;

  i_i_8 <= i_i_3 + const_expression_2;

  
  out0_102 <= '1' WHEN i_i_8 > to_unsigned(16#10#, 8) ELSE
      '0';

  
  j_j_8 <= j_j_3 WHEN out0_102 = '0' ELSE
      j_j_4;

  
  out0_86 <= '1' WHEN j_j_8 > to_unsigned(16#20#, 8) ELSE
      '0';

  
  sit_30 <= sit_20 WHEN out0_86 = '0' ELSE
      sit_1;

  
  out0_1 <= '1' WHEN sit_20 = to_unsigned(16#0C#, 8) ELSE
      '0';

  
  out0_118 <= sit WHEN out0_1 = '0' ELSE
      sit_30;

  
  out0_3 <= '1' WHEN sit_20 = to_unsigned(16#0B#, 8) ELSE
      '0';

  
  out0_119 <= out0_118 WHEN out0_3 = '0' ELSE
      sit_2;

  
  out0_5 <= '1' WHEN sit_20 = to_unsigned(16#0A#, 8) ELSE
      '0';

  
  out0_120 <= out0_119 WHEN out0_5 = '0' ELSE
      sit_29;

  
  out0_7 <= '1' WHEN sit_20 = to_unsigned(16#09#, 8) ELSE
      '0';

  
  out0_121 <= out0_120 WHEN out0_7 = '0' ELSE
      sit_28;

  
  out0_9 <= '1' WHEN sit_20 = to_unsigned(16#08#, 8) ELSE
      '0';

  
  out0_122 <= out0_121 WHEN out0_9 = '0' ELSE
      sit_27;

  
  out0_11 <= '1' WHEN sit_20 = to_unsigned(16#06#, 8) ELSE
      '0';

  
  out0_123 <= out0_122 WHEN out0_11 = '0' ELSE
      sit_26;

  
  out0_13 <= '1' WHEN sit_20 = to_unsigned(16#05#, 8) ELSE
      '0';

  
  out0_124 <= out0_123 WHEN out0_13 = '0' ELSE
      sit_9;

  
  out0_15 <= '1' WHEN sit_20 = to_unsigned(16#04#, 8) ELSE
      '0';

  
  out0_125 <= out0_124 WHEN out0_15 = '0' ELSE
      sit_25;

  
  out0_17 <= '1' WHEN sit_20 = to_unsigned(16#27#, 8) ELSE
      '0';

  
  out0_126 <= out0_125 WHEN out0_17 = '0' ELSE
      sit_12;

  
  out0_19 <= '1' WHEN sit_20 = to_unsigned(16#20#, 8) ELSE
      '0';

  
  out0_127 <= out0_126 WHEN out0_19 = '0' ELSE
      sit_24;

  
  out0_21 <= '1' WHEN sit_20 = to_unsigned(16#1F#, 8) ELSE
      '0';

  
  out0_128 <= out0_127 WHEN out0_21 = '0' ELSE
      sit_14;

  
  out0_23 <= '1' WHEN sit_20 = to_unsigned(16#03#, 8) ELSE
      '0';

  
  out0_129 <= out0_128 WHEN out0_23 = '0' ELSE
      sit_15;

  
  out0_25 <= '1' WHEN sit_20 = to_unsigned(16#15#, 8) ELSE
      '0';

  
  out0_130 <= out0_129 WHEN out0_25 = '0' ELSE
      sit_16;

  
  out0_27 <= '1' WHEN sit_20 = to_unsigned(16#02#, 8) ELSE
      '0';

  
  out0_131 <= out0_130 WHEN out0_27 = '0' ELSE
      sit_17;

  
  out0_29 <= '1' WHEN sit_20 = to_unsigned(16#01#, 8) ELSE
      '0';

  
  out0_132 <= out0_131 WHEN out0_29 = '0' ELSE
      sit_23;

  
  sit_out <= out0_132 WHEN out0_31 = '0' ELSE
      sit_22;

  intdelay6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        sit_20 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        sit_20 <= sit_out;
      END IF;
    END IF;
  END PROCESS intdelay6_process;


  -- %
  
  out0_31 <= '1' WHEN sit_20 = to_unsigned(16#00#, 8) ELSE
      '0';

  valid_out_1 <= '0';

  valid_out_2 <= '1';

  
  out0_133 <= valid_out_1 WHEN out0_1 = '0' ELSE
      valid_out_2;

  valid_out_3 <= '0';

  
  out0_134 <= out0_133 WHEN out0_3 = '0' ELSE
      valid_out_3;

  valid_out_4 <= '0';

  
  out0_135 <= out0_134 WHEN out0_5 = '0' ELSE
      valid_out_4;

  valid_out_5 <= '0';

  
  out0_136 <= out0_135 WHEN out0_7 = '0' ELSE
      valid_out_5;

  valid_out_6 <= '0';

  
  out0_137 <= out0_136 WHEN out0_9 = '0' ELSE
      valid_out_6;

  valid_out_7 <= '0';

  
  out0_138 <= out0_137 WHEN out0_11 = '0' ELSE
      valid_out_7;

  valid_out_8 <= '0';

  
  out0_139 <= out0_138 WHEN out0_13 = '0' ELSE
      valid_out_8;

  valid_out_9 <= '0';

  
  out0_140 <= out0_139 WHEN out0_15 = '0' ELSE
      valid_out_9;

  valid_out_10 <= '0';

  
  out0_141 <= out0_140 WHEN out0_17 = '0' ELSE
      valid_out_10;

  valid_out_11 <= '0';

  
  out0_142 <= out0_141 WHEN out0_19 = '0' ELSE
      valid_out_11;

  valid_out_12 <= '0';

  
  out0_143 <= out0_142 WHEN out0_21 = '0' ELSE
      valid_out_12;

  valid_out_13 <= '0';

  
  out0_144 <= out0_143 WHEN out0_23 = '0' ELSE
      valid_out_13;

  valid_out_14 <= '0';

  
  out0_145 <= out0_144 WHEN out0_25 = '0' ELSE
      valid_out_14;

  valid_out_15 <= '0';

  
  out0_146 <= out0_145 WHEN out0_27 = '0' ELSE
      valid_out_15;

  valid_out_16 <= '0';

  
  out0_147 <= out0_146 WHEN out0_29 = '0' ELSE
      valid_out_16;

  valid_out_17 <= '0';

  
  valid_out_18 <= out0_147 WHEN out0_31 = '0' ELSE
      valid_out_17;

  Unit_Delay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Unit_Delay4_out1 <= '0';
      ELSIF enb = '1' THEN
        Unit_Delay4_out1 <= valid_out_18;
      END IF;
    END IF;
  END PROCESS Unit_Delay4_process;


  
  Data_Type_Conversion_out1 <= '1' WHEN Unit_Delay4_out1 /= '0' ELSE
      '0';

  valid_out <= Data_Type_Conversion_out1;

  data_out_re <= X"00000000";
  data_out_im <= X"00000000";

  ram_out_re <= X"00000000";
  ram_out_im <= X"00000000";

  ram_out_re_1 <= X"00000000";
  ram_out_im_1 <= X"00000000";

  
  out0_re <= ram_out_re WHEN out0_1 = '0' ELSE
      ram_out_re_1;
  
  out0_im <= ram_out_im WHEN out0_1 = '0' ELSE
      ram_out_im_1;

  ram_out_re_2 <= X"00000000";
  ram_out_im_2 <= X"00000000";

  
  out0_re_1 <= out0_re WHEN out0_3 = '0' ELSE
      ram_out_re_2;
  
  out0_im_1 <= out0_im WHEN out0_3 = '0' ELSE
      ram_out_im_2;

  ram_out_re_3 <= X"00000000";
  ram_out_im_3 <= X"00000000";

  
  out0_re_2 <= out0_re_1 WHEN out0_5 = '0' ELSE
      ram_out_re_3;
  
  out0_im_2 <= out0_im_1 WHEN out0_5 = '0' ELSE
      ram_out_im_3;

  ram_out_re_4 <= X"00000000";
  ram_out_im_4 <= X"00000000";

  
  out0_re_3 <= out0_re_2 WHEN out0_7 = '0' ELSE
      ram_out_re_4;
  
  out0_im_3 <= out0_im_2 WHEN out0_7 = '0' ELSE
      ram_out_im_4;

  
  relop1_relop1 <= '1' WHEN i_i_3 /= j_j_3 ELSE
      '0';

  ram_out_re_5 <= X"00000000";
  ram_out_im_5 <= X"00000000";

  
  relop_relop1 <= '1' WHEN i_i_3 /= j_j_3 ELSE
      '0';

  ram_out_re_6 <= X"00000000";
  ram_out_im_6 <= X"00000000";

  ram_out_re_7 <= X"00000000";
  ram_out_im_7 <= X"00000000";

  ram_out_re_8 <= X"00000000";
  ram_out_im_8 <= X"00000000";

  ram_out_re_9 <= X"00000000";
  ram_out_im_9 <= X"00000000";

  ram_out_re_10 <= X"00000000";
  ram_out_im_10 <= X"00000000";

  ram_out_re_11 <= X"00000000";
  ram_out_im_11 <= X"00000000";

  ram_out_re_12 <= X"00000000";
  ram_out_im_12 <= X"00000000";

  ram_out_re_13 <= X"00000000";
  ram_out_im_13 <= X"00000000";

  ram_out_re_14 <= X"3f800000";
  ram_out_im_14 <= X"00000000";

  ram_out_re_15 <= X"00000000";
  ram_out_im_15 <= X"00000000";

  Unit_Delay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Unit_Delay3_out1_re <= X"00000000";
        Unit_Delay3_out1_im <= X"00000000";
      ELSIF enb = '1' THEN
        Unit_Delay3_out1_re <= in_ri_re;
        Unit_Delay3_out1_im <= in_ri_im;
      END IF;
    END IF;
  END PROCESS Unit_Delay3_process;


  
  ram_out_re_16 <= ram_out_re_15 WHEN out0 = '0' ELSE
      Unit_Delay3_out1_re;
  
  ram_out_im_16 <= ram_out_im_15 WHEN out0 = '0' ELSE
      Unit_Delay3_out1_im;

  we <= '0';

  we_1 <= '0';

  
  out0_148 <= we WHEN out0_1 = '0' ELSE
      we_1;

  we_2 <= '0';

  
  out0_149 <= out0_148 WHEN out0_3 = '0' ELSE
      we_2;

  we_3 <= '0';

  
  out0_150 <= out0_149 WHEN out0_5 = '0' ELSE
      we_3;

  we_4 <= '0';

  
  out0_151 <= out0_150 WHEN out0_7 = '0' ELSE
      we_4;

  we_5 <= '0';

  we_6 <= '1';

  
  we_7 <= we_5 WHEN relop1_relop1 = '0' ELSE
      we_6;

  
  out0_152 <= out0_151 WHEN out0_9 = '0' ELSE
      we_7;

  we_8 <= '0';

  
  out0_153 <= out0_152 WHEN out0_11 = '0' ELSE
      we_8;

  we_9 <= '0';

  
  out0_154 <= out0_153 WHEN out0_13 = '0' ELSE
      we_9;

  we_10 <= '0';

  
  out0_155 <= out0_154 WHEN out0_15 = '0' ELSE
      we_10;

  we_11 <= '1';

  
  out0_156 <= out0_155 WHEN out0_17 = '0' ELSE
      we_11;

  we_12 <= '0';

  
  out0_157 <= out0_156 WHEN out0_19 = '0' ELSE
      we_12;

  we_13 <= '0';

  
  out0_158 <= out0_157 WHEN out0_21 = '0' ELSE
      we_13;

  we_14 <= '0';

  
  out0_159 <= out0_158 WHEN out0_23 = '0' ELSE
      we_14;

  we_15 <= '0';

  
  out0_160 <= out0_159 WHEN out0_25 = '0' ELSE
      we_15;

  we_16 <= '0';

  
  out0_161 <= out0_160 WHEN out0_27 = '0' ELSE
      we_16;

  we_17 <= '1';

  
  out0_162 <= out0_161 WHEN out0_29 = '0' ELSE
      we_17;

  we_18 <= '0';

  we_19 <= '1';

  
  we_20 <= we_18 WHEN out0 = '0' ELSE
      we_19;

  
  we_21 <= out0_162 WHEN out0_31 = '0' ELSE
      we_20;

  ram_add1 <= to_unsigned(16#0000#, 16);

  j_j_11 <= resize(j_j_9, 16);

  jj <= j_j_11 sll 4;

  i_i_11 <= resize(i_i_9, 16);

  ram_add1_1 <= jj + i_i_11;

  
  out0_163 <= ram_add1 WHEN out0_1 = '0' ELSE
      ram_add1_1;

  j_j_12 <= resize(j_j_3, 16);

  jj_1 <= j_j_12 sll 4;

  i_i_12 <= resize(i_i_3, 16);

  ram_add1_2 <= jj_1 + i_i_12;

  
  out0_164 <= out0_163 WHEN out0_3 = '0' ELSE
      ram_add1_2;

  ram_add1_3 <= to_unsigned(16#0000#, 16);

  
  out0_165 <= out0_164 WHEN out0_5 = '0' ELSE
      ram_add1_3;

  ram_add1_4 <= to_unsigned(16#0000#, 16);

  
  out0_166 <= out0_165 WHEN out0_7 = '0' ELSE
      ram_add1_4;

  ram_add1_5 <= to_unsigned(16#0000#, 16);

  j_j_13 <= resize(k_k_3, 16);

  jj_2 <= j_j_13 sll 4;

  i_i_13 <= resize(j_j_3, 16);

  ram_add1_6 <= jj_2 + i_i_13;

  
  ram_add1_7 <= ram_add1_5 WHEN relop1_relop1 = '0' ELSE
      ram_add1_6;

  
  out0_167 <= out0_166 WHEN out0_9 = '0' ELSE
      ram_add1_7;

  j_j_14 <= resize(i_i_3, 16);

  jj_3 <= j_j_14 sll 4;

  i_i_14 <= resize(j_j_3, 16);

  ram_add1_8 <= jj_3 + i_i_14;

  
  out0_168 <= out0_167 WHEN out0_11 = '0' ELSE
      ram_add1_8;

  j_j_15 <= resize(i_i_3, 16);

  jj_4 <= j_j_15 sll 4;

  i_i_15 <= resize(j_j_3, 16);

  ram_add1_9 <= jj_4 + i_i_15;

  
  out0_169 <= out0_168 WHEN out0_13 = '0' ELSE
      ram_add1_9;

  ram_add1_10 <= to_unsigned(16#0000#, 16);

  
  out0_170 <= out0_169 WHEN out0_15 = '0' ELSE
      ram_add1_10;

  j_j_16 <= resize(k_k_3, 16);

  jj_5 <= j_j_16 sll 4;

  i_i_16 <= resize(i_i_3, 16);

  ram_add1_11 <= jj_5 + i_i_16;

  
  out0_171 <= out0_170 WHEN out0_17 = '0' ELSE
      ram_add1_11;

  ram_add1_12 <= to_unsigned(16#0000#, 16);

  
  out0_172 <= out0_171 WHEN out0_19 = '0' ELSE
      ram_add1_12;

  ram_add1_13 <= to_unsigned(16#0000#, 16);

  
  out0_173 <= out0_172 WHEN out0_21 = '0' ELSE
      ram_add1_13;

  j_j_17 <= resize(k_k_3, 16);

  jj_6 <= j_j_17 sll 4;

  i_i_17 <= resize(i_i_3, 16);

  ram_add1_14 <= jj_6 + i_i_17;

  
  out0_174 <= out0_173 WHEN out0_23 = '0' ELSE
      ram_add1_14;

  ram_add1_15 <= to_unsigned(16#0000#, 16);

  
  out0_175 <= out0_174 WHEN out0_25 = '0' ELSE
      ram_add1_15;

  j_j_18 <= resize(i_i_3, 16);

  jj_7 <= j_j_18 sll 4;

  i_i_18 <= resize(i_i_3, 16);

  ram_add1_16 <= jj_7 + i_i_18;

  
  out0_176 <= out0_175 WHEN out0_27 = '0' ELSE
      ram_add1_16;

  n_n <= to_unsigned(16#10#, 8);

  out0_177 <= n_n + i_i_3;

  j_j_19 <= resize(out0_177, 16);

  jj_8 <= j_j_19 sll 4;

  i_i_19 <= resize(i_i_3, 16);

  ram_add1_17 <= jj_8 + i_i_19;

  
  out0_178 <= out0_176 WHEN out0_29 = '0' ELSE
      ram_add1_17;

  ram_add1_18 <= to_unsigned(16#0000#, 16);

  j_j_20 <= resize(j1, 16);

  jj_9 <= j_j_20 sll 4;

  i_i_20 <= resize(i1_3, 16);

  ram_add1_19 <= jj_9 + i_i_20;

  
  ram_add1_20 <= ram_add1_18 WHEN out0 = '0' ELSE
      ram_add1_19;

  
  ram_add1_21 <= out0_178 WHEN out0_31 = '0' ELSE
      ram_add1_20;

  ram_add2 <= to_unsigned(16#0000#, 16);

  j_j_21 <= resize(j_j_9, 16);

  jj_10 <= j_j_21 sll 4;

  i_i_21 <= resize(i_i_9, 16);

  ram_add2_1 <= jj_10 + i_i_21;

  
  out0_179 <= ram_add2 WHEN out0_1 = '0' ELSE
      ram_add2_1;

  j_j_22 <= resize(j_j_3, 16);

  jj_11 <= j_j_22 sll 4;

  i_i_22 <= resize(i_i_3, 16);

  ram_add2_2 <= jj_11 + i_i_22;

  
  out0_180 <= out0_179 WHEN out0_3 = '0' ELSE
      ram_add2_2;

  ram_add2_3 <= to_unsigned(16#0000#, 16);

  
  out0_181 <= out0_180 WHEN out0_5 = '0' ELSE
      ram_add2_3;

  ram_add2_4 <= to_unsigned(16#0000#, 16);

  
  out0_182 <= out0_181 WHEN out0_7 = '0' ELSE
      ram_add2_4;

  ram_add2_5 <= to_unsigned(16#0000#, 16);

  j_j_23 <= resize(k_k_3, 16);

  jj_12 <= j_j_23 sll 4;

  i_i_23 <= resize(j_j_3, 16);

  ram_add2_6 <= jj_12 + i_i_23;

  
  ram_add2_7 <= ram_add2_5 WHEN relop1_relop1 = '0' ELSE
      ram_add2_6;

  
  out0_183 <= out0_182 WHEN out0_9 = '0' ELSE
      ram_add2_7;

  j_j_24 <= resize(k_k_7, 16);

  jj_13 <= j_j_24 sll 4;

  i_i_24 <= resize(i_i_3, 16);

  ram_add2_8 <= jj_13 + i_i_24;

  
  out0_184 <= out0_183 WHEN out0_11 = '0' ELSE
      ram_add2_8;

  j_j_25 <= resize(k_k_3, 16);

  jj_14 <= j_j_25 sll 4;

  i_i_25 <= resize(i_i_3, 16);

  ram_add2_9 <= jj_14 + i_i_25;

  
  out0_185 <= out0_184 WHEN out0_13 = '0' ELSE
      ram_add2_9;

  ram_add2_10 <= to_unsigned(16#0000#, 16);

  
  out0_186 <= out0_185 WHEN out0_15 = '0' ELSE
      ram_add2_10;

  j_j_26 <= resize(k_k_3, 16);

  jj_15 <= j_j_26 sll 4;

  i_i_26 <= resize(i_i_3, 16);

  ram_add2_11 <= jj_15 + i_i_26;

  
  out0_187 <= out0_186 WHEN out0_17 = '0' ELSE
      ram_add2_11;

  ram_add2_12 <= to_unsigned(16#0000#, 16);

  
  out0_188 <= out0_187 WHEN out0_19 = '0' ELSE
      ram_add2_12;

  ram_add2_13 <= to_unsigned(16#0000#, 16);

  
  out0_189 <= out0_188 WHEN out0_21 = '0' ELSE
      ram_add2_13;

  j_j_27 <= resize(k_k_3, 16);

  jj_16 <= j_j_27 sll 4;

  i_i_27 <= resize(i_i_3, 16);

  ram_add2_14 <= jj_16 + i_i_27;

  
  out0_190 <= out0_189 WHEN out0_23 = '0' ELSE
      ram_add2_14;

  ram_add2_15 <= to_unsigned(16#0000#, 16);

  
  out0_191 <= out0_190 WHEN out0_25 = '0' ELSE
      ram_add2_15;

  j_j_28 <= resize(i_i_3, 16);

  jj_17 <= j_j_28 sll 4;

  i_i_28 <= resize(i_i_3, 16);

  ram_add2_16 <= jj_17 + i_i_28;

  
  out0_192 <= out0_191 WHEN out0_27 = '0' ELSE
      ram_add2_16;

  n_n_1 <= to_unsigned(16#10#, 8);

  out0_193 <= n_n_1 + i_i_3;

  j_j_29 <= resize(out0_193, 16);

  jj_18 <= j_j_29 sll 4;

  i_i_29 <= resize(i_i_3, 16);

  ram_add2_17 <= jj_18 + i_i_29;

  
  out0_194 <= out0_192 WHEN out0_29 = '0' ELSE
      ram_add2_17;

  ram_add2_18 <= to_unsigned(16#0000#, 16);

  j_j_30 <= resize(j1, 16);

  jj_19 <= j_j_30 sll 4;

  i_i_30 <= resize(i1_3, 16);

  ram_add2_19 <= jj_19 + i_i_30;

  
  ram_add2_20 <= ram_add2_18 WHEN out0 = '0' ELSE
      ram_add2_19;

  
  ram_add2_21 <= out0_194 WHEN out0_31 = '0' ELSE
      ram_add2_20;

  ram_add3 <= to_unsigned(16#0000#, 16);

  j_j_31 <= resize(j_j_9, 16);

  jj_20 <= j_j_31 sll 4;

  i_i_31 <= resize(i_i_9, 16);

  ram_add3_1 <= jj_20 + i_i_31;

  
  out0_195 <= ram_add3 WHEN out0_1 = '0' ELSE
      ram_add3_1;

  j_j_32 <= resize(j_j_3, 16);

  jj_21 <= j_j_32 sll 4;

  i_i_32 <= resize(i_i_3, 16);

  ram_add3_2 <= jj_21 + i_i_32;

  
  out0_196 <= out0_195 WHEN out0_3 = '0' ELSE
      ram_add3_2;

  ram_add3_3 <= to_unsigned(16#0000#, 16);

  
  out0_197 <= out0_196 WHEN out0_5 = '0' ELSE
      ram_add3_3;

  ram_add3_4 <= to_unsigned(16#0000#, 16);

  
  out0_198 <= out0_197 WHEN out0_7 = '0' ELSE
      ram_add3_4;

  ram_add3_5 <= to_unsigned(16#0000#, 16);

  j_j_33 <= resize(k_k_3, 16);

  jj_22 <= j_j_33 sll 4;

  i_i_33 <= resize(j_j_3, 16);

  ram_add3_6 <= jj_22 + i_i_33;

  
  ram_add3_7 <= ram_add3_5 WHEN relop1_relop1 = '0' ELSE
      ram_add3_6;

  
  out0_199 <= out0_198 WHEN out0_9 = '0' ELSE
      ram_add3_7;

  j_j_34 <= resize(k_k_7, 16);

  jj_23 <= j_j_34 sll 4;

  i_i_34 <= resize(j_j_3, 16);

  ram_add3_8 <= jj_23 + i_i_34;

  
  out0_200 <= out0_199 WHEN out0_11 = '0' ELSE
      ram_add3_8;

  j_j_35 <= resize(k_k_3, 16);

  jj_24 <= j_j_35 sll 4;

  i_i_35 <= resize(j_j_3, 16);

  ram_add3_9 <= jj_24 + i_i_35;

  
  out0_201 <= out0_200 WHEN out0_13 = '0' ELSE
      ram_add3_9;

  ram_add3_10 <= to_unsigned(16#0000#, 16);

  
  out0_202 <= out0_201 WHEN out0_15 = '0' ELSE
      ram_add3_10;

  j_j_36 <= resize(k_k_3, 16);

  jj_25 <= j_j_36 sll 4;

  i_i_36 <= resize(i_i_3, 16);

  ram_add3_11 <= jj_25 + i_i_36;

  
  out0_203 <= out0_202 WHEN out0_17 = '0' ELSE
      ram_add3_11;

  ram_add3_12 <= to_unsigned(16#0000#, 16);

  
  out0_204 <= out0_203 WHEN out0_19 = '0' ELSE
      ram_add3_12;

  ram_add3_13 <= to_unsigned(16#0000#, 16);

  
  out0_205 <= out0_204 WHEN out0_21 = '0' ELSE
      ram_add3_13;

  j_j_37 <= resize(k_k_3, 16);

  jj_26 <= j_j_37 sll 4;

  i_i_37 <= resize(i_i_3, 16);

  ram_add3_14 <= jj_26 + i_i_37;

  
  out0_206 <= out0_205 WHEN out0_23 = '0' ELSE
      ram_add3_14;

  ram_add3_15 <= to_unsigned(16#0000#, 16);

  
  out0_207 <= out0_206 WHEN out0_25 = '0' ELSE
      ram_add3_15;

  j_j_38 <= resize(i_i_3, 16);

  jj_27 <= j_j_38 sll 4;

  i_i_38 <= resize(i_i_3, 16);

  ram_add3_16 <= jj_27 + i_i_38;

  
  out0_208 <= out0_207 WHEN out0_27 = '0' ELSE
      ram_add3_16;

  n_n_2 <= to_unsigned(16#10#, 8);

  out0_209 <= n_n_2 + i_i_3;

  j_j_39 <= resize(out0_209, 16);

  jj_28 <= j_j_39 sll 4;

  i_i_39 <= resize(i_i_3, 16);

  ram_add3_17 <= jj_28 + i_i_39;

  
  out0_210 <= out0_208 WHEN out0_29 = '0' ELSE
      ram_add3_17;

  ram_add3_18 <= to_unsigned(16#0000#, 16);

  j_j_40 <= resize(j1, 16);

  jj_29 <= j_j_40 sll 4;

  i_i_40 <= resize(i1_3, 16);

  ram_add3_19 <= jj_29 + i_i_40;

  
  ram_add3_20 <= ram_add3_18 WHEN out0 = '0' ELSE
      ram_add3_19;

  
  ram_add3_21 <= out0_210 WHEN out0_31 = '0' ELSE
      ram_add3_20;

  intdelay10_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        p2_re <= X"00000000";
        p2_im <= X"00000000";
      ELSIF enb = '1' THEN
        p2_re <= dout2_re;
        p2_im <= dout2_im;
      END IF;
    END IF;
  END PROCESS intdelay10_process;


  
  out0_re_4 <= p2_re WHEN out0_1 = '0' ELSE
      p2_re;
  
  out0_im_4 <= p2_im WHEN out0_1 = '0' ELSE
      p2_im;

  
  out0_re_5 <= out0_re_4 WHEN out0_3 = '0' ELSE
      p2_re;
  
  out0_im_5 <= out0_im_4 WHEN out0_3 = '0' ELSE
      p2_im;

  
  out0_re_6 <= out0_re_5 WHEN out0_5 = '0' ELSE
      p2_re;
  
  out0_im_6 <= out0_im_5 WHEN out0_5 = '0' ELSE
      p2_im;

  
  out0_re_7 <= out0_re_6 WHEN out0_7 = '0' ELSE
      p2_re;
  
  out0_im_7 <= out0_im_6 WHEN out0_7 = '0' ELSE
      p2_im;

  
  out0_re_8 <= out0_re_7 WHEN out0_9 = '0' ELSE
      p2_re;
  
  out0_im_8 <= out0_im_7 WHEN out0_9 = '0' ELSE
      p2_im;

  
  out0_re_9 <= out0_re_8 WHEN out0_11 = '0' ELSE
      p2_re;
  
  out0_im_9 <= out0_im_8 WHEN out0_11 = '0' ELSE
      p2_im;

  
  out0_re_10 <= out0_re_9 WHEN out0_13 = '0' ELSE
      p2_re;
  
  out0_im_10 <= out0_im_9 WHEN out0_13 = '0' ELSE
      p2_im;

  
  out0_re_11 <= out0_re_10 WHEN out0_15 = '0' ELSE
      p2_re;
  
  out0_im_11 <= out0_im_10 WHEN out0_15 = '0' ELSE
      p2_im;

  
  out0_re_12 <= out0_re_11 WHEN out0_17 = '0' ELSE
      p2_re;
  
  out0_im_12 <= out0_im_11 WHEN out0_17 = '0' ELSE
      p2_im;

  
  out0_re_13 <= out0_re_12 WHEN out0_19 = '0' ELSE
      p2_re;
  
  out0_im_13 <= out0_im_12 WHEN out0_19 = '0' ELSE
      p2_im;

  
  out0_re_14 <= out0_re_13 WHEN out0_21 = '0' ELSE
      memory_out1_re;
  
  out0_im_14 <= out0_im_13 WHEN out0_21 = '0' ELSE
      memory_out1_im;

  
  out0_re_15 <= out0_re_14 WHEN out0_23 = '0' ELSE
      p2_re;
  
  out0_im_15 <= out0_im_14 WHEN out0_23 = '0' ELSE
      p2_im;

  
  out0_re_16 <= out0_re_15 WHEN out0_25 = '0' ELSE
      p2_re;
  
  out0_im_16 <= out0_im_15 WHEN out0_25 = '0' ELSE
      p2_im;

  
  out0_re_17 <= out0_re_16 WHEN out0_27 = '0' ELSE
      p2_re;
  
  out0_im_17 <= out0_im_16 WHEN out0_27 = '0' ELSE
      p2_im;

  
  out0_re_18 <= out0_re_17 WHEN out0_29 = '0' ELSE
      p2_re;
  
  out0_im_18 <= out0_im_17 WHEN out0_29 = '0' ELSE
      p2_im;

  
  dout2_re <= out0_re_18 WHEN out0_31 = '0' ELSE
      p2_re;
  
  dout2_im <= out0_im_18 WHEN out0_31 = '0' ELSE
      p2_im;

  -- #codegen
  intdelay11_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        p1_re <= X"00000000";
        p1_im <= X"00000000";
      ELSIF enb = '1' THEN
        p1_re <= dout1_re;
        p1_im <= dout1_im;
      END IF;
    END IF;
  END PROCESS intdelay11_process;


  
  out0_re_19 <= p1_re WHEN out0_1 = '0' ELSE
      p1_re;
  
  out0_im_19 <= p1_im WHEN out0_1 = '0' ELSE
      p1_im;

  
  out0_re_20 <= out0_re_19 WHEN out0_3 = '0' ELSE
      p1_re;
  
  out0_im_20 <= out0_im_19 WHEN out0_3 = '0' ELSE
      p1_im;

  
  out0_re_21 <= out0_re_20 WHEN out0_5 = '0' ELSE
      p1_re;
  
  out0_im_21 <= out0_im_20 WHEN out0_5 = '0' ELSE
      p1_im;

  
  out0_re_22 <= out0_re_21 WHEN out0_7 = '0' ELSE
      p1_re;
  
  out0_im_22 <= out0_im_21 WHEN out0_7 = '0' ELSE
      p1_im;

  
  out0_re_23 <= out0_re_22 WHEN out0_9 = '0' ELSE
      p1_re;
  
  out0_im_23 <= out0_im_22 WHEN out0_9 = '0' ELSE
      p1_im;

  
  out0_re_24 <= out0_re_23 WHEN out0_11 = '0' ELSE
      p1_re;
  
  out0_im_24 <= out0_im_23 WHEN out0_11 = '0' ELSE
      p1_im;

  
  out0_re_25 <= out0_re_24 WHEN out0_13 = '0' ELSE
      p1_re;
  
  out0_im_25 <= out0_im_24 WHEN out0_13 = '0' ELSE
      p1_im;

  
  out0_re_26 <= out0_re_25 WHEN out0_15 = '0' ELSE
      p1_re;
  
  out0_im_26 <= out0_im_25 WHEN out0_15 = '0' ELSE
      p1_im;

  
  out0_re_27 <= out0_re_26 WHEN out0_17 = '0' ELSE
      p1_re;
  
  out0_im_27 <= out0_im_26 WHEN out0_17 = '0' ELSE
      p1_im;

  
  out0_re_28 <= out0_re_27 WHEN out0_19 = '0' ELSE
      p1_re;
  
  out0_im_28 <= out0_im_27 WHEN out0_19 = '0' ELSE
      p1_im;

  
  out0_re_29 <= out0_re_28 WHEN out0_21 = '0' ELSE
      p1_re;
  
  out0_im_29 <= out0_im_28 WHEN out0_21 = '0' ELSE
      p1_im;

  
  out0_re_30 <= out0_re_29 WHEN out0_23 = '0' ELSE
      p1_re;
  
  out0_im_30 <= out0_im_29 WHEN out0_23 = '0' ELSE
      p1_im;

  
  out0_re_31 <= out0_re_30 WHEN out0_25 = '0' ELSE
      memory_out1_re;
  
  out0_im_31 <= out0_im_30 WHEN out0_25 = '0' ELSE
      memory_out1_im;

  
  out0_re_32 <= out0_re_31 WHEN out0_27 = '0' ELSE
      p1_re;
  
  out0_im_32 <= out0_im_31 WHEN out0_27 = '0' ELSE
      p1_im;

  
  out0_re_33 <= out0_re_32 WHEN out0_29 = '0' ELSE
      p1_re;
  
  out0_im_33 <= out0_im_32 WHEN out0_29 = '0' ELSE
      p1_im;

  
  dout1_re <= out0_re_33 WHEN out0_31 = '0' ELSE
      p1_re;
  
  dout1_im <= out0_im_33 WHEN out0_31 = '0' ELSE
      p1_im;

  
  p5_re_1 <= p5_re WHEN relop_relop1 = '0' ELSE
      memory_out3_re;
  
  p5_im_1 <= p5_im WHEN relop_relop1 = '0' ELSE
      memory_out3_im;

  intdelay7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        p5_re <= X"00000000";
        p5_im <= X"00000000";
      ELSIF enb = '1' THEN
        p5_re <= dout5_re;
        p5_im <= dout5_im;
      END IF;
    END IF;
  END PROCESS intdelay7_process;


  
  out0_re_34 <= p5_re WHEN out0_1 = '0' ELSE
      p5_re;
  
  out0_im_34 <= p5_im WHEN out0_1 = '0' ELSE
      p5_im;

  
  out0_re_35 <= out0_re_34 WHEN out0_3 = '0' ELSE
      p5_re;
  
  out0_im_35 <= out0_im_34 WHEN out0_3 = '0' ELSE
      p5_im;

  
  out0_re_36 <= out0_re_35 WHEN out0_5 = '0' ELSE
      p5_re;
  
  out0_im_36 <= out0_im_35 WHEN out0_5 = '0' ELSE
      p5_im;

  
  out0_re_37 <= out0_re_36 WHEN out0_7 = '0' ELSE
      p5_re;
  
  out0_im_37 <= out0_im_36 WHEN out0_7 = '0' ELSE
      p5_im;

  
  out0_re_38 <= out0_re_37 WHEN out0_9 = '0' ELSE
      p5_re;
  
  out0_im_38 <= out0_im_37 WHEN out0_9 = '0' ELSE
      p5_im;

  
  out0_re_39 <= out0_re_38 WHEN out0_11 = '0' ELSE
      p5_re_1;
  
  out0_im_39 <= out0_im_38 WHEN out0_11 = '0' ELSE
      p5_im_1;

  
  out0_re_40 <= out0_re_39 WHEN out0_13 = '0' ELSE
      p5_re;
  
  out0_im_40 <= out0_im_39 WHEN out0_13 = '0' ELSE
      p5_im;

  
  out0_re_41 <= out0_re_40 WHEN out0_15 = '0' ELSE
      p5_re;
  
  out0_im_41 <= out0_im_40 WHEN out0_15 = '0' ELSE
      p5_im;

  
  out0_re_42 <= out0_re_41 WHEN out0_17 = '0' ELSE
      p5_re;
  
  out0_im_42 <= out0_im_41 WHEN out0_17 = '0' ELSE
      p5_im;

  
  out0_re_43 <= out0_re_42 WHEN out0_19 = '0' ELSE
      p5_re;
  
  out0_im_43 <= out0_im_42 WHEN out0_19 = '0' ELSE
      p5_im;

  
  out0_re_44 <= out0_re_43 WHEN out0_21 = '0' ELSE
      p5_re;
  
  out0_im_44 <= out0_im_43 WHEN out0_21 = '0' ELSE
      p5_im;

  
  out0_re_45 <= out0_re_44 WHEN out0_23 = '0' ELSE
      p5_re;
  
  out0_im_45 <= out0_im_44 WHEN out0_23 = '0' ELSE
      p5_im;

  
  out0_re_46 <= out0_re_45 WHEN out0_25 = '0' ELSE
      p5_re;
  
  out0_im_46 <= out0_im_45 WHEN out0_25 = '0' ELSE
      p5_im;

  
  out0_re_47 <= out0_re_46 WHEN out0_27 = '0' ELSE
      p5_re;
  
  out0_im_47 <= out0_im_46 WHEN out0_27 = '0' ELSE
      p5_im;

  
  out0_re_48 <= out0_re_47 WHEN out0_29 = '0' ELSE
      p5_re;
  
  out0_im_48 <= out0_im_47 WHEN out0_29 = '0' ELSE
      p5_im;

  
  dout5_re <= out0_re_48 WHEN out0_31 = '0' ELSE
      p5_re;
  
  dout5_im <= out0_im_48 WHEN out0_31 = '0' ELSE
      p5_im;

  
  p4_re_1 <= p4_re WHEN relop_relop1 = '0' ELSE
      memory_out2_re;
  
  p4_im_1 <= p4_im WHEN relop_relop1 = '0' ELSE
      memory_out2_im;

  intdelay8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        p4_re <= X"00000000";
        p4_im <= X"00000000";
      ELSIF enb = '1' THEN
        p4_re <= dout4_re;
        p4_im <= dout4_im;
      END IF;
    END IF;
  END PROCESS intdelay8_process;


  
  out0_re_49 <= p4_re WHEN out0_1 = '0' ELSE
      p4_re;
  
  out0_im_49 <= p4_im WHEN out0_1 = '0' ELSE
      p4_im;

  
  out0_re_50 <= out0_re_49 WHEN out0_3 = '0' ELSE
      p4_re;
  
  out0_im_50 <= out0_im_49 WHEN out0_3 = '0' ELSE
      p4_im;

  
  out0_re_51 <= out0_re_50 WHEN out0_5 = '0' ELSE
      p4_re;
  
  out0_im_51 <= out0_im_50 WHEN out0_5 = '0' ELSE
      p4_im;

  
  out0_re_52 <= out0_re_51 WHEN out0_7 = '0' ELSE
      p4_re;
  
  out0_im_52 <= out0_im_51 WHEN out0_7 = '0' ELSE
      p4_im;

  
  out0_re_53 <= out0_re_52 WHEN out0_9 = '0' ELSE
      p4_re;
  
  out0_im_53 <= out0_im_52 WHEN out0_9 = '0' ELSE
      p4_im;

  
  out0_re_54 <= out0_re_53 WHEN out0_11 = '0' ELSE
      p4_re_1;
  
  out0_im_54 <= out0_im_53 WHEN out0_11 = '0' ELSE
      p4_im_1;

  
  out0_re_55 <= out0_re_54 WHEN out0_13 = '0' ELSE
      p4_re;
  
  out0_im_55 <= out0_im_54 WHEN out0_13 = '0' ELSE
      p4_im;

  
  out0_re_56 <= out0_re_55 WHEN out0_15 = '0' ELSE
      p4_re;
  
  out0_im_56 <= out0_im_55 WHEN out0_15 = '0' ELSE
      p4_im;

  
  out0_re_57 <= out0_re_56 WHEN out0_17 = '0' ELSE
      p4_re;
  
  out0_im_57 <= out0_im_56 WHEN out0_17 = '0' ELSE
      p4_im;

  
  out0_re_58 <= out0_re_57 WHEN out0_19 = '0' ELSE
      p4_re;
  
  out0_im_58 <= out0_im_57 WHEN out0_19 = '0' ELSE
      p4_im;

  
  out0_re_59 <= out0_re_58 WHEN out0_21 = '0' ELSE
      p4_re;
  
  out0_im_59 <= out0_im_58 WHEN out0_21 = '0' ELSE
      p4_im;

  
  out0_re_60 <= out0_re_59 WHEN out0_23 = '0' ELSE
      p4_re;
  
  out0_im_60 <= out0_im_59 WHEN out0_23 = '0' ELSE
      p4_im;

  
  out0_re_61 <= out0_re_60 WHEN out0_25 = '0' ELSE
      p4_re;
  
  out0_im_61 <= out0_im_60 WHEN out0_25 = '0' ELSE
      p4_im;

  
  out0_re_62 <= out0_re_61 WHEN out0_27 = '0' ELSE
      p4_re;
  
  out0_im_62 <= out0_im_61 WHEN out0_27 = '0' ELSE
      p4_im;

  
  out0_re_63 <= out0_re_62 WHEN out0_29 = '0' ELSE
      p4_re;
  
  out0_im_63 <= out0_im_62 WHEN out0_29 = '0' ELSE
      p4_im;

  
  dout4_re <= out0_re_63 WHEN out0_31 = '0' ELSE
      p4_re;
  
  dout4_im <= out0_im_63 WHEN out0_31 = '0' ELSE
      p4_im;

  
  p3_re_1 <= p3_re WHEN relop_relop1 = '0' ELSE
      memory_out1_re;
  
  p3_im_1 <= p3_im WHEN relop_relop1 = '0' ELSE
      memory_out1_im;

  intdelay9_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        p3_re <= X"00000000";
        p3_im <= X"00000000";
      ELSIF enb = '1' THEN
        p3_re <= dout3_re;
        p3_im <= dout3_im;
      END IF;
    END IF;
  END PROCESS intdelay9_process;


  
  out0_re_64 <= p3_re WHEN out0_1 = '0' ELSE
      p3_re;
  
  out0_im_64 <= p3_im WHEN out0_1 = '0' ELSE
      p3_im;

  
  out0_re_65 <= out0_re_64 WHEN out0_3 = '0' ELSE
      p3_re;
  
  out0_im_65 <= out0_im_64 WHEN out0_3 = '0' ELSE
      p3_im;

  
  out0_re_66 <= out0_re_65 WHEN out0_5 = '0' ELSE
      p3_re;
  
  out0_im_66 <= out0_im_65 WHEN out0_5 = '0' ELSE
      p3_im;

  
  out0_re_67 <= out0_re_66 WHEN out0_7 = '0' ELSE
      p3_re;
  
  out0_im_67 <= out0_im_66 WHEN out0_7 = '0' ELSE
      p3_im;

  
  out0_re_68 <= out0_re_67 WHEN out0_9 = '0' ELSE
      p3_re;
  
  out0_im_68 <= out0_im_67 WHEN out0_9 = '0' ELSE
      p3_im;

  
  out0_re_69 <= out0_re_68 WHEN out0_11 = '0' ELSE
      p3_re_1;
  
  out0_im_69 <= out0_im_68 WHEN out0_11 = '0' ELSE
      p3_im_1;

  
  out0_re_70 <= out0_re_69 WHEN out0_13 = '0' ELSE
      p3_re;
  
  out0_im_70 <= out0_im_69 WHEN out0_13 = '0' ELSE
      p3_im;

  
  out0_re_71 <= out0_re_70 WHEN out0_15 = '0' ELSE
      p3_re;
  
  out0_im_71 <= out0_im_70 WHEN out0_15 = '0' ELSE
      p3_im;

  
  out0_re_72 <= out0_re_71 WHEN out0_17 = '0' ELSE
      p3_re;
  
  out0_im_72 <= out0_im_71 WHEN out0_17 = '0' ELSE
      p3_im;

  
  out0_re_73 <= out0_re_72 WHEN out0_19 = '0' ELSE
      p3_re;
  
  out0_im_73 <= out0_im_72 WHEN out0_19 = '0' ELSE
      p3_im;

  
  out0_re_74 <= out0_re_73 WHEN out0_21 = '0' ELSE
      p3_re;
  
  out0_im_74 <= out0_im_73 WHEN out0_21 = '0' ELSE
      p3_im;

  
  out0_re_75 <= out0_re_74 WHEN out0_23 = '0' ELSE
      p3_re;
  
  out0_im_75 <= out0_im_74 WHEN out0_23 = '0' ELSE
      p3_im;

  
  out0_re_76 <= out0_re_75 WHEN out0_25 = '0' ELSE
      p3_re;
  
  out0_im_76 <= out0_im_75 WHEN out0_25 = '0' ELSE
      p3_im;

  
  out0_re_77 <= out0_re_76 WHEN out0_27 = '0' ELSE
      p3_re;
  
  out0_im_77 <= out0_im_76 WHEN out0_27 = '0' ELSE
      p3_im;

  
  out0_re_78 <= out0_re_77 WHEN out0_29 = '0' ELSE
      p3_re;
  
  out0_im_78 <= out0_im_77 WHEN out0_29 = '0' ELSE
      p3_im;

  
  dout3_re <= out0_re_78 WHEN out0_31 = '0' ELSE
      p3_re;
  
  dout3_im <= out0_im_78 WHEN out0_31 = '0' ELSE
      p3_im;

  
  ram_out_re_17 <= ram_out_re_5 WHEN relop1_relop1 = '0' ELSE
      func2_out1_re;
  
  ram_out_im_17 <= ram_out_im_5 WHEN relop1_relop1 = '0' ELSE
      func2_out1_im;

  
  out0_re_79 <= out0_re_3 WHEN out0_9 = '0' ELSE
      ram_out_re_17;
  
  out0_im_79 <= out0_im_3 WHEN out0_9 = '0' ELSE
      ram_out_im_17;

  
  out0_re_80 <= out0_re_79 WHEN out0_11 = '0' ELSE
      ram_out_re_6;
  
  out0_im_80 <= out0_im_79 WHEN out0_11 = '0' ELSE
      ram_out_im_6;

  
  out0_re_81 <= out0_re_80 WHEN out0_13 = '0' ELSE
      ram_out_re_7;
  
  out0_im_81 <= out0_im_80 WHEN out0_13 = '0' ELSE
      ram_out_im_7;

  
  out0_re_82 <= out0_re_81 WHEN out0_15 = '0' ELSE
      ram_out_re_8;
  
  out0_im_82 <= out0_im_81 WHEN out0_15 = '0' ELSE
      ram_out_im_8;

  
  out0_re_83 <= out0_re_82 WHEN out0_17 = '0' ELSE
      func1_out1_re;
  
  out0_im_83 <= out0_im_82 WHEN out0_17 = '0' ELSE
      func1_out1_im;

  
  out0_re_84 <= out0_re_83 WHEN out0_19 = '0' ELSE
      ram_out_re_9;
  
  out0_im_84 <= out0_im_83 WHEN out0_19 = '0' ELSE
      ram_out_im_9;

  
  out0_re_85 <= out0_re_84 WHEN out0_21 = '0' ELSE
      ram_out_re_10;
  
  out0_im_85 <= out0_im_84 WHEN out0_21 = '0' ELSE
      ram_out_im_10;

  
  out0_re_86 <= out0_re_85 WHEN out0_23 = '0' ELSE
      ram_out_re_11;
  
  out0_im_86 <= out0_im_85 WHEN out0_23 = '0' ELSE
      ram_out_im_11;

  
  out0_re_87 <= out0_re_86 WHEN out0_25 = '0' ELSE
      ram_out_re_12;
  
  out0_im_87 <= out0_im_86 WHEN out0_25 = '0' ELSE
      ram_out_im_12;

  
  out0_re_88 <= out0_re_87 WHEN out0_27 = '0' ELSE
      ram_out_re_13;
  
  out0_im_88 <= out0_im_87 WHEN out0_27 = '0' ELSE
      ram_out_im_13;

  
  out0_re_89 <= out0_re_88 WHEN out0_29 = '0' ELSE
      ram_out_re_14;
  
  out0_im_89 <= out0_im_88 WHEN out0_29 = '0' ELSE
      ram_out_im_14;

  
  ram_out_re_18 <= out0_re_89 WHEN out0_31 = '0' ELSE
      ram_out_re_16;
  
  ram_out_im_18 <= out0_im_89 WHEN out0_31 = '0' ELSE
      ram_out_im_16;

  
  out0_re_90 <= data_out_re WHEN out0_1 = '0' ELSE
      memory_out1_re;
  
  out0_im_90 <= data_out_im WHEN out0_1 = '0' ELSE
      memory_out1_im;

  data_out_re_1 <= X"00000000";
  data_out_im_1 <= X"00000000";

  
  out0_re_91 <= out0_re_90 WHEN out0_3 = '0' ELSE
      data_out_re_1;
  
  out0_im_91 <= out0_im_90 WHEN out0_3 = '0' ELSE
      data_out_im_1;

  data_out_re_2 <= X"00000000";
  data_out_im_2 <= X"00000000";

  
  out0_re_92 <= out0_re_91 WHEN out0_5 = '0' ELSE
      data_out_re_2;
  
  out0_im_92 <= out0_im_91 WHEN out0_5 = '0' ELSE
      data_out_im_2;

  data_out_re_3 <= X"00000000";
  data_out_im_3 <= X"00000000";

  
  out0_re_93 <= out0_re_92 WHEN out0_7 = '0' ELSE
      data_out_re_3;
  
  out0_im_93 <= out0_im_92 WHEN out0_7 = '0' ELSE
      data_out_im_3;

  data_out_re_4 <= X"00000000";
  data_out_im_4 <= X"00000000";

  
  out0_re_94 <= out0_re_93 WHEN out0_9 = '0' ELSE
      data_out_re_4;
  
  out0_im_94 <= out0_im_93 WHEN out0_9 = '0' ELSE
      data_out_im_4;

  data_out_re_5 <= X"00000000";
  data_out_im_5 <= X"00000000";

  
  out0_re_95 <= out0_re_94 WHEN out0_11 = '0' ELSE
      data_out_re_5;
  
  out0_im_95 <= out0_im_94 WHEN out0_11 = '0' ELSE
      data_out_im_5;

  data_out_re_6 <= X"00000000";
  data_out_im_6 <= X"00000000";

  
  out0_re_96 <= out0_re_95 WHEN out0_13 = '0' ELSE
      data_out_re_6;
  
  out0_im_96 <= out0_im_95 WHEN out0_13 = '0' ELSE
      data_out_im_6;

  data_out_re_7 <= X"00000000";
  data_out_im_7 <= X"00000000";

  
  out0_re_97 <= out0_re_96 WHEN out0_15 = '0' ELSE
      data_out_re_7;
  
  out0_im_97 <= out0_im_96 WHEN out0_15 = '0' ELSE
      data_out_im_7;

  data_out_re_8 <= X"00000000";
  data_out_im_8 <= X"00000000";

  
  out0_re_98 <= out0_re_97 WHEN out0_17 = '0' ELSE
      data_out_re_8;
  
  out0_im_98 <= out0_im_97 WHEN out0_17 = '0' ELSE
      data_out_im_8;

  data_out_re_9 <= X"00000000";
  data_out_im_9 <= X"00000000";

  
  out0_re_99 <= out0_re_98 WHEN out0_19 = '0' ELSE
      data_out_re_9;
  
  out0_im_99 <= out0_im_98 WHEN out0_19 = '0' ELSE
      data_out_im_9;

  data_out_re_10 <= X"00000000";
  data_out_im_10 <= X"00000000";

  
  out0_re_100 <= out0_re_99 WHEN out0_21 = '0' ELSE
      data_out_re_10;
  
  out0_im_100 <= out0_im_99 WHEN out0_21 = '0' ELSE
      data_out_im_10;

  data_out_re_11 <= X"00000000";
  data_out_im_11 <= X"00000000";

  
  out0_re_101 <= out0_re_100 WHEN out0_23 = '0' ELSE
      data_out_re_11;
  
  out0_im_101 <= out0_im_100 WHEN out0_23 = '0' ELSE
      data_out_im_11;

  data_out_re_12 <= X"00000000";
  data_out_im_12 <= X"00000000";

  
  out0_re_102 <= out0_re_101 WHEN out0_25 = '0' ELSE
      data_out_re_12;
  
  out0_im_102 <= out0_im_101 WHEN out0_25 = '0' ELSE
      data_out_im_12;

  data_out_re_13 <= X"00000000";
  data_out_im_13 <= X"00000000";

  
  out0_re_103 <= out0_re_102 WHEN out0_27 = '0' ELSE
      data_out_re_13;
  
  out0_im_103 <= out0_im_102 WHEN out0_27 = '0' ELSE
      data_out_im_13;

  data_out_re_14 <= X"00000000";
  data_out_im_14 <= X"00000000";

  
  out0_re_104 <= out0_re_103 WHEN out0_29 = '0' ELSE
      data_out_re_14;
  
  out0_im_104 <= out0_im_103 WHEN out0_29 = '0' ELSE
      data_out_im_14;

  data_out_re_15 <= X"00000000";
  data_out_im_15 <= X"00000000";

  
  data_out_re_16 <= out0_re_104 WHEN out0_31 = '0' ELSE
      data_out_re_15;
  
  data_out_im_16 <= out0_im_104 WHEN out0_31 = '0' ELSE
      data_out_im_15;

  Unit_Delay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Unit_Delay1_out1_re <= X"00000000";
        Unit_Delay1_out1_im <= X"00000000";
      ELSIF enb = '1' THEN
        Unit_Delay1_out1_re <= data_out_re_16;
        Unit_Delay1_out1_im <= data_out_im_16;
      END IF;
    END IF;
  END PROCESS Unit_Delay1_process;


  ce_out <= clk_enable;

  out_ir_re <= Unit_Delay1_out1_re;

  out_ir_im <= Unit_Delay1_out1_im;

END rtl;

