LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY SimpleDualPortRAM_generic IS
  GENERIC( AddrWidth                      : integer := 1;
           DataWidth                      : integer := 1
           );
  PORT( clk                               :   IN    std_logic;
        wr_din                            :   IN    std_logic_vector(DataWidth - 1 DOWNTO 0);
        wr_addr                           :   IN    std_logic_vector(AddrWidth - 1 DOWNTO 0);
        wr_en                             :   IN    std_logic;
        rd_addr                           :   IN    std_logic_vector(AddrWidth - 1 DOWNTO 0);
        rd_dout                           :   OUT   std_logic_vector(DataWidth - 1 DOWNTO 0)
        );
END SimpleDualPortRAM_generic;


ARCHITECTURE rtl OF SimpleDualPortRAM_generic IS

  -- Local Type Definitions
  TYPE ram_type IS ARRAY (2**AddrWidth - 1 DOWNTO 0) of std_logic_vector(DataWidth - 1 DOWNTO 0);

  -- Signals
  SIGNAL ram                              : ram_type;
  SIGNAL data_int                         : std_logic_vector(DataWidth - 1 DOWNTO 0);
  SIGNAL wr_addr_unsigned                 : unsigned(AddrWidth - 1 DOWNTO 0);
  SIGNAL rd_addr_unsigned                 : unsigned(AddrWidth - 1 DOWNTO 0);

BEGIN
  wr_addr_unsigned <= unsigned(wr_addr);

  rd_addr_unsigned <= unsigned(rd_addr);

  ShiftRegisterRAM_Wrapper_generic_process: PROCESS (clk)
  BEGIN
    IF clk'event AND clk = '1' THEN
      IF wr_en = '1' THEN
        ram(to_integer(wr_addr_unsigned)) <= wr_din;
      END IF;
      data_int <= ram(to_integer(rd_addr_unsigned));
    END IF;
  END PROCESS ShiftRegisterRAM_Wrapper_generic_process;

  rd_dout <= data_int;

END rtl;

